magic
tech sky130A
magscale 1 2
timestamp 1718283729
<< metal3 >>
rect -1186 1012 1248 1040
rect -1186 -1012 1164 1012
rect 1228 -1012 1248 1012
rect -1186 -1040 1248 -1012
<< via3 >>
rect 1164 -1012 1228 1012
<< mimcap >>
rect -1146 960 854 1000
rect -1146 -960 -1106 960
rect 814 -960 854 960
rect -1146 -1000 854 -960
<< mimcapcontact >>
rect -1106 -960 814 960
<< metal4 >>
rect 1148 1012 1244 1028
rect -1107 960 815 961
rect -1107 -960 -1106 960
rect 814 -960 815 960
rect -1107 -961 815 -960
rect 1148 -1012 1164 1012
rect 1228 -1012 1244 1012
rect 1148 -1028 1244 -1012
<< properties >>
string FIXED_BBOX -1186 -1040 894 1040
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10.00 l 10.00 val 207.6 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
