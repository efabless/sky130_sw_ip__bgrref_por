magic
tech sky130A
magscale 1 2
timestamp 1718283729
<< error_p >>
rect -29 138 29 144
rect -29 104 -17 138
rect -29 98 29 104
rect -29 -104 29 -98
rect -29 -138 -17 -104
rect -29 -144 29 -138
<< pwell >>
rect -211 -260 211 260
<< nmos >>
rect -15 -50 15 50
<< ndiff >>
rect -73 38 -15 50
rect -73 -38 -61 38
rect -27 -38 -15 38
rect -73 -50 -15 -38
rect 15 38 73 50
rect 15 -38 27 38
rect 61 -38 73 38
rect 15 -50 73 -38
<< ndiffc >>
rect -61 -38 -27 38
rect 27 -38 61 38
<< psubdiff >>
rect -175 190 -79 224
rect 79 190 175 224
rect -175 128 -141 190
rect 141 128 175 190
rect -175 -190 -141 -128
rect 141 -190 175 -128
rect -175 -224 -79 -190
rect 79 -224 175 -190
<< psubdiffcont >>
rect -79 190 79 224
rect -175 -128 -141 128
rect 141 -128 175 128
rect -79 -224 79 -190
<< poly >>
rect -33 138 33 154
rect -33 104 -17 138
rect 17 104 33 138
rect -33 88 33 104
rect -15 50 15 88
rect -15 -88 15 -50
rect -33 -104 33 -88
rect -33 -138 -17 -104
rect 17 -138 33 -104
rect -33 -154 33 -138
<< polycont >>
rect -17 104 17 138
rect -17 -138 17 -104
<< locali >>
rect -175 190 -79 224
rect 79 190 175 224
rect -175 128 -141 190
rect -33 104 -17 138
rect 17 104 33 138
rect 141 128 175 190
rect -61 38 -27 54
rect -61 -54 -27 -38
rect 27 38 61 54
rect 27 -54 61 -38
rect -175 -190 -141 -128
rect -33 -138 -17 -104
rect 17 -138 33 -104
rect 141 -190 175 -128
rect -175 -224 -79 -190
rect 79 -224 175 -190
<< viali >>
rect -17 104 17 138
rect -61 -38 -27 38
rect 27 -38 61 38
rect -17 -138 17 -104
<< metal1 >>
rect -29 138 29 144
rect -29 104 -17 138
rect 17 104 29 138
rect -29 98 29 104
rect -67 38 -21 50
rect -67 -38 -61 38
rect -27 -38 -21 38
rect -67 -50 -21 -38
rect 21 38 67 50
rect 21 -38 27 38
rect 61 -38 67 38
rect 21 -50 67 -38
rect -29 -104 29 -98
rect -29 -138 -17 -104
rect 17 -138 29 -104
rect -29 -144 29 -138
<< properties >>
string FIXED_BBOX -158 -207 158 207
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
