magic
tech sky130A
magscale 1 2
timestamp 1717527227
<< pwell >>
rect -1363 -1582 1363 1582
<< psubdiff >>
rect -1327 1512 -1231 1546
rect 1231 1512 1327 1546
rect -1327 1450 -1293 1512
rect 1293 1450 1327 1512
rect -1327 -1512 -1293 -1450
rect 1293 -1512 1327 -1450
rect -1327 -1546 -1231 -1512
rect 1231 -1546 1327 -1512
<< psubdiffcont >>
rect -1231 1512 1231 1546
rect -1327 -1450 -1293 1450
rect 1293 -1450 1327 1450
rect -1231 -1546 1231 -1512
<< xpolycontact >>
rect -1197 984 -1127 1416
rect -1197 -1416 -1127 -984
rect -1031 984 -961 1416
rect -1031 -1416 -961 -984
rect -865 984 -795 1416
rect -865 -1416 -795 -984
rect -699 984 -629 1416
rect -699 -1416 -629 -984
rect -533 984 -463 1416
rect -533 -1416 -463 -984
rect -367 984 -297 1416
rect -367 -1416 -297 -984
rect -201 984 -131 1416
rect -201 -1416 -131 -984
rect -35 984 35 1416
rect -35 -1416 35 -984
rect 131 984 201 1416
rect 131 -1416 201 -984
rect 297 984 367 1416
rect 297 -1416 367 -984
rect 463 984 533 1416
rect 463 -1416 533 -984
rect 629 984 699 1416
rect 629 -1416 699 -984
rect 795 984 865 1416
rect 795 -1416 865 -984
rect 961 984 1031 1416
rect 961 -1416 1031 -984
rect 1127 984 1197 1416
rect 1127 -1416 1197 -984
<< xpolyres >>
rect -1197 -984 -1127 984
rect -1031 -984 -961 984
rect -865 -984 -795 984
rect -699 -984 -629 984
rect -533 -984 -463 984
rect -367 -984 -297 984
rect -201 -984 -131 984
rect -35 -984 35 984
rect 131 -984 201 984
rect 297 -984 367 984
rect 463 -984 533 984
rect 629 -984 699 984
rect 795 -984 865 984
rect 961 -984 1031 984
rect 1127 -984 1197 984
<< locali >>
rect -1327 1512 -1231 1546
rect 1231 1512 1327 1546
rect -1327 1450 -1293 1512
rect 1293 1450 1327 1512
rect -1327 -1512 -1293 -1450
rect 1293 -1512 1327 -1450
rect -1327 -1546 -1231 -1512
rect 1231 -1546 1327 -1512
<< viali >>
rect -1181 1001 -1143 1398
rect -1015 1001 -977 1398
rect -849 1001 -811 1398
rect -683 1001 -645 1398
rect -517 1001 -479 1398
rect -351 1001 -313 1398
rect -185 1001 -147 1398
rect -19 1001 19 1398
rect 147 1001 185 1398
rect 313 1001 351 1398
rect 479 1001 517 1398
rect 645 1001 683 1398
rect 811 1001 849 1398
rect 977 1001 1015 1398
rect 1143 1001 1181 1398
rect -1181 -1398 -1143 -1001
rect -1015 -1398 -977 -1001
rect -849 -1398 -811 -1001
rect -683 -1398 -645 -1001
rect -517 -1398 -479 -1001
rect -351 -1398 -313 -1001
rect -185 -1398 -147 -1001
rect -19 -1398 19 -1001
rect 147 -1398 185 -1001
rect 313 -1398 351 -1001
rect 479 -1398 517 -1001
rect 645 -1398 683 -1001
rect 811 -1398 849 -1001
rect 977 -1398 1015 -1001
rect 1143 -1398 1181 -1001
<< metal1 >>
rect -1187 1398 -1137 1410
rect -1187 1001 -1181 1398
rect -1143 1001 -1137 1398
rect -1187 989 -1137 1001
rect -1021 1398 -971 1410
rect -1021 1001 -1015 1398
rect -977 1001 -971 1398
rect -1021 989 -971 1001
rect -855 1398 -805 1410
rect -855 1001 -849 1398
rect -811 1001 -805 1398
rect -855 989 -805 1001
rect -689 1398 -639 1410
rect -689 1001 -683 1398
rect -645 1001 -639 1398
rect -689 989 -639 1001
rect -523 1398 -473 1410
rect -523 1001 -517 1398
rect -479 1001 -473 1398
rect -523 989 -473 1001
rect -357 1398 -307 1410
rect -357 1001 -351 1398
rect -313 1001 -307 1398
rect -357 989 -307 1001
rect -191 1398 -141 1410
rect -191 1001 -185 1398
rect -147 1001 -141 1398
rect -191 989 -141 1001
rect -25 1398 25 1410
rect -25 1001 -19 1398
rect 19 1001 25 1398
rect -25 989 25 1001
rect 141 1398 191 1410
rect 141 1001 147 1398
rect 185 1001 191 1398
rect 141 989 191 1001
rect 307 1398 357 1410
rect 307 1001 313 1398
rect 351 1001 357 1398
rect 307 989 357 1001
rect 473 1398 523 1410
rect 473 1001 479 1398
rect 517 1001 523 1398
rect 473 989 523 1001
rect 639 1398 689 1410
rect 639 1001 645 1398
rect 683 1001 689 1398
rect 639 989 689 1001
rect 805 1398 855 1410
rect 805 1001 811 1398
rect 849 1001 855 1398
rect 805 989 855 1001
rect 971 1398 1021 1410
rect 971 1001 977 1398
rect 1015 1001 1021 1398
rect 971 989 1021 1001
rect 1137 1398 1187 1410
rect 1137 1001 1143 1398
rect 1181 1001 1187 1398
rect 1137 989 1187 1001
rect -1187 -1001 -1137 -989
rect -1187 -1398 -1181 -1001
rect -1143 -1398 -1137 -1001
rect -1187 -1410 -1137 -1398
rect -1021 -1001 -971 -989
rect -1021 -1398 -1015 -1001
rect -977 -1398 -971 -1001
rect -1021 -1410 -971 -1398
rect -855 -1001 -805 -989
rect -855 -1398 -849 -1001
rect -811 -1398 -805 -1001
rect -855 -1410 -805 -1398
rect -689 -1001 -639 -989
rect -689 -1398 -683 -1001
rect -645 -1398 -639 -1001
rect -689 -1410 -639 -1398
rect -523 -1001 -473 -989
rect -523 -1398 -517 -1001
rect -479 -1398 -473 -1001
rect -523 -1410 -473 -1398
rect -357 -1001 -307 -989
rect -357 -1398 -351 -1001
rect -313 -1398 -307 -1001
rect -357 -1410 -307 -1398
rect -191 -1001 -141 -989
rect -191 -1398 -185 -1001
rect -147 -1398 -141 -1001
rect -191 -1410 -141 -1398
rect -25 -1001 25 -989
rect -25 -1398 -19 -1001
rect 19 -1398 25 -1001
rect -25 -1410 25 -1398
rect 141 -1001 191 -989
rect 141 -1398 147 -1001
rect 185 -1398 191 -1001
rect 141 -1410 191 -1398
rect 307 -1001 357 -989
rect 307 -1398 313 -1001
rect 351 -1398 357 -1001
rect 307 -1410 357 -1398
rect 473 -1001 523 -989
rect 473 -1398 479 -1001
rect 517 -1398 523 -1001
rect 473 -1410 523 -1398
rect 639 -1001 689 -989
rect 639 -1398 645 -1001
rect 683 -1398 689 -1001
rect 639 -1410 689 -1398
rect 805 -1001 855 -989
rect 805 -1398 811 -1001
rect 849 -1398 855 -1001
rect 805 -1410 855 -1398
rect 971 -1001 1021 -989
rect 971 -1398 977 -1001
rect 1015 -1398 1021 -1001
rect 971 -1410 1021 -1398
rect 1137 -1001 1187 -989
rect 1137 -1398 1143 -1001
rect 1181 -1398 1187 -1001
rect 1137 -1410 1187 -1398
<< properties >>
string FIXED_BBOX -1310 -1529 1310 1529
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 10.0 m 1 nx 15 wmin 0.350 lmin 0.50 rho 2000 val 58.218k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
