magic
tech sky130A
magscale 1 2
timestamp 1717363523
<< pwell >>
rect -201 -15582 201 15582
<< psubdiff >>
rect -165 15512 -69 15546
rect 69 15512 165 15546
rect -165 15450 -131 15512
rect 131 15450 165 15512
rect -165 -15512 -131 -15450
rect 131 -15512 165 -15450
rect -165 -15546 -69 -15512
rect 69 -15546 165 -15512
<< psubdiffcont >>
rect -69 15512 69 15546
rect -165 -15450 -131 15450
rect 131 -15450 165 15450
rect -69 -15546 69 -15512
<< xpolycontact >>
rect -35 14984 35 15416
rect -35 -15416 35 -14984
<< xpolyres >>
rect -35 -14984 35 14984
<< locali >>
rect -165 15512 -69 15546
rect 69 15512 165 15546
rect -165 15450 -131 15512
rect 131 15450 165 15512
rect -165 -15512 -131 -15450
rect 131 -15512 165 -15450
rect -165 -15546 -69 -15512
rect 69 -15546 165 -15512
<< viali >>
rect -19 15001 19 15398
rect -19 -15398 19 -15001
<< metal1 >>
rect -25 15398 25 15410
rect -25 15001 -19 15398
rect 19 15001 25 15398
rect -25 14989 25 15001
rect -25 -15001 25 -14989
rect -25 -15398 -19 -15001
rect 19 -15398 25 -15001
rect -25 -15410 25 -15398
<< properties >>
string FIXED_BBOX -148 -15529 148 15529
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 150.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 858.218k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
