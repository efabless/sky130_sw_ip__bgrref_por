magic
tech sky130A
magscale 1 2
timestamp 1717527227
<< error_p >>
rect -1295 122 -1237 128
rect -1295 88 -1283 122
rect -1295 82 -1237 88
<< pwell >>
rect -1463 -260 1463 260
<< nmos >>
rect -1263 -50 -1233 50
rect -1167 -50 -1137 50
rect -1071 -50 -1041 50
rect -975 -50 -945 50
rect -879 -50 -849 50
rect -783 -50 -753 50
rect -687 -50 -657 50
rect -591 -50 -561 50
rect -495 -50 -465 50
rect -399 -50 -369 50
rect -303 -50 -273 50
rect -207 -50 -177 50
rect -111 -50 -81 50
rect -15 -50 15 50
rect 81 -50 111 50
rect 177 -50 207 50
rect 273 -50 303 50
rect 369 -50 399 50
rect 465 -50 495 50
rect 561 -50 591 50
rect 657 -50 687 50
rect 753 -50 783 50
rect 849 -50 879 50
rect 945 -50 975 50
rect 1041 -50 1071 50
rect 1137 -50 1167 50
rect 1233 -50 1263 50
<< ndiff >>
rect -1325 38 -1263 50
rect -1325 -38 -1313 38
rect -1279 -38 -1263 38
rect -1325 -50 -1263 -38
rect -1233 38 -1167 50
rect -1233 -38 -1217 38
rect -1183 -38 -1167 38
rect -1233 -50 -1167 -38
rect -1137 38 -1071 50
rect -1137 -38 -1121 38
rect -1087 -38 -1071 38
rect -1137 -50 -1071 -38
rect -1041 38 -975 50
rect -1041 -38 -1025 38
rect -991 -38 -975 38
rect -1041 -50 -975 -38
rect -945 38 -879 50
rect -945 -38 -929 38
rect -895 -38 -879 38
rect -945 -50 -879 -38
rect -849 38 -783 50
rect -849 -38 -833 38
rect -799 -38 -783 38
rect -849 -50 -783 -38
rect -753 38 -687 50
rect -753 -38 -737 38
rect -703 -38 -687 38
rect -753 -50 -687 -38
rect -657 38 -591 50
rect -657 -38 -641 38
rect -607 -38 -591 38
rect -657 -50 -591 -38
rect -561 38 -495 50
rect -561 -38 -545 38
rect -511 -38 -495 38
rect -561 -50 -495 -38
rect -465 38 -399 50
rect -465 -38 -449 38
rect -415 -38 -399 38
rect -465 -50 -399 -38
rect -369 38 -303 50
rect -369 -38 -353 38
rect -319 -38 -303 38
rect -369 -50 -303 -38
rect -273 38 -207 50
rect -273 -38 -257 38
rect -223 -38 -207 38
rect -273 -50 -207 -38
rect -177 38 -111 50
rect -177 -38 -161 38
rect -127 -38 -111 38
rect -177 -50 -111 -38
rect -81 38 -15 50
rect -81 -38 -65 38
rect -31 -38 -15 38
rect -81 -50 -15 -38
rect 15 38 81 50
rect 15 -38 31 38
rect 65 -38 81 38
rect 15 -50 81 -38
rect 111 38 177 50
rect 111 -38 127 38
rect 161 -38 177 38
rect 111 -50 177 -38
rect 207 38 273 50
rect 207 -38 223 38
rect 257 -38 273 38
rect 207 -50 273 -38
rect 303 38 369 50
rect 303 -38 319 38
rect 353 -38 369 38
rect 303 -50 369 -38
rect 399 38 465 50
rect 399 -38 415 38
rect 449 -38 465 38
rect 399 -50 465 -38
rect 495 38 561 50
rect 495 -38 511 38
rect 545 -38 561 38
rect 495 -50 561 -38
rect 591 38 657 50
rect 591 -38 607 38
rect 641 -38 657 38
rect 591 -50 657 -38
rect 687 38 753 50
rect 687 -38 703 38
rect 737 -38 753 38
rect 687 -50 753 -38
rect 783 38 849 50
rect 783 -38 799 38
rect 833 -38 849 38
rect 783 -50 849 -38
rect 879 38 945 50
rect 879 -38 895 38
rect 929 -38 945 38
rect 879 -50 945 -38
rect 975 38 1041 50
rect 975 -38 991 38
rect 1025 -38 1041 38
rect 975 -50 1041 -38
rect 1071 38 1137 50
rect 1071 -38 1087 38
rect 1121 -38 1137 38
rect 1071 -50 1137 -38
rect 1167 38 1233 50
rect 1167 -38 1183 38
rect 1217 -38 1233 38
rect 1167 -50 1233 -38
rect 1263 38 1325 50
rect 1263 -38 1279 38
rect 1313 -38 1325 38
rect 1263 -50 1325 -38
<< ndiffc >>
rect -1313 -38 -1279 38
rect -1217 -38 -1183 38
rect -1121 -38 -1087 38
rect -1025 -38 -991 38
rect -929 -38 -895 38
rect -833 -38 -799 38
rect -737 -38 -703 38
rect -641 -38 -607 38
rect -545 -38 -511 38
rect -449 -38 -415 38
rect -353 -38 -319 38
rect -257 -38 -223 38
rect -161 -38 -127 38
rect -65 -38 -31 38
rect 31 -38 65 38
rect 127 -38 161 38
rect 223 -38 257 38
rect 319 -38 353 38
rect 415 -38 449 38
rect 511 -38 545 38
rect 607 -38 641 38
rect 703 -38 737 38
rect 799 -38 833 38
rect 895 -38 929 38
rect 991 -38 1025 38
rect 1087 -38 1121 38
rect 1183 -38 1217 38
rect 1279 -38 1313 38
<< psubdiff >>
rect -1427 190 -1331 224
rect 1331 190 1427 224
rect -1427 128 -1393 190
rect 1393 128 1427 190
rect -1427 -190 -1393 -128
rect 1393 -190 1427 -128
rect -1427 -224 -1331 -190
rect 1331 -224 1427 -190
<< psubdiffcont >>
rect -1331 190 1331 224
rect -1427 -128 -1393 128
rect 1393 -128 1427 128
rect -1331 -224 1331 -190
<< poly >>
rect -1299 122 -1233 138
rect -1299 88 -1283 122
rect -1249 88 -1233 122
rect -1299 72 -1233 88
rect -1263 50 -1233 72
rect -1167 122 -1041 138
rect -1167 88 -1150 122
rect -1057 88 -1041 122
rect -1167 72 -1041 88
rect -1167 50 -1137 72
rect -1071 50 -1041 72
rect -975 122 -273 138
rect -975 88 -949 122
rect -299 88 -273 122
rect -975 72 -273 88
rect -975 50 -945 72
rect -879 50 -849 72
rect -783 50 -753 72
rect -687 50 -657 72
rect -591 50 -561 72
rect -495 50 -465 72
rect -399 50 -369 72
rect -303 50 -273 72
rect -207 122 1263 138
rect -207 88 -181 122
rect 1237 88 1263 122
rect -207 72 1263 88
rect -207 50 -177 72
rect -111 50 -81 72
rect -15 50 15 72
rect 81 50 111 72
rect 177 50 207 72
rect 273 50 303 72
rect 369 50 399 72
rect 465 50 495 72
rect 561 50 591 72
rect 657 50 687 72
rect 753 50 783 72
rect 849 50 879 72
rect 945 50 975 72
rect 1041 50 1071 72
rect 1137 50 1167 72
rect 1233 50 1263 72
rect -1263 -76 -1233 -50
rect -1167 -76 -1137 -50
rect -1071 -76 -1041 -50
rect -975 -76 -945 -50
rect -879 -76 -849 -50
rect -783 -76 -753 -50
rect -687 -76 -657 -50
rect -591 -76 -561 -50
rect -495 -76 -465 -50
rect -399 -76 -369 -50
rect -303 -76 -273 -50
rect -207 -76 -177 -50
rect -111 -76 -81 -50
rect -15 -76 15 -50
rect 81 -76 111 -50
rect 177 -76 207 -50
rect 273 -76 303 -50
rect 369 -76 399 -50
rect 465 -76 495 -50
rect 561 -76 591 -50
rect 657 -76 687 -50
rect 753 -76 783 -50
rect 849 -76 879 -50
rect 945 -76 975 -50
rect 1041 -76 1071 -50
rect 1137 -76 1167 -50
rect 1233 -76 1263 -50
<< polycont >>
rect -1283 88 -1249 122
rect -1150 88 -1057 122
rect -949 88 -299 122
rect -181 88 1237 122
<< locali >>
rect -1427 190 -1331 224
rect 1331 190 1427 224
rect -1427 128 -1393 190
rect 1393 128 1427 190
rect -1299 88 -1283 122
rect -1249 88 -1233 122
rect -1167 88 -1150 122
rect -1057 88 -1041 122
rect -975 88 -949 122
rect -299 88 -273 122
rect -207 88 -181 122
rect 1237 88 1263 122
rect -1313 38 -1279 54
rect -1313 -54 -1279 -38
rect -1217 38 -1183 54
rect -1217 -54 -1183 -38
rect -1121 38 -1087 54
rect -1121 -54 -1087 -38
rect -1025 38 -991 54
rect -1025 -54 -991 -38
rect -929 38 -895 54
rect -929 -54 -895 -38
rect -833 38 -799 54
rect -833 -54 -799 -38
rect -737 38 -703 54
rect -737 -54 -703 -38
rect -641 38 -607 54
rect -641 -54 -607 -38
rect -545 38 -511 54
rect -545 -54 -511 -38
rect -449 38 -415 54
rect -449 -54 -415 -38
rect -353 38 -319 54
rect -353 -54 -319 -38
rect -257 38 -223 54
rect -257 -54 -223 -38
rect -161 38 -127 54
rect -161 -54 -127 -38
rect -65 38 -31 54
rect -65 -54 -31 -38
rect 31 38 65 54
rect 31 -54 65 -38
rect 127 38 161 54
rect 127 -54 161 -38
rect 223 38 257 54
rect 223 -54 257 -38
rect 319 38 353 54
rect 319 -54 353 -38
rect 415 38 449 54
rect 415 -54 449 -38
rect 511 38 545 54
rect 511 -54 545 -38
rect 607 38 641 54
rect 607 -54 641 -38
rect 703 38 737 54
rect 703 -54 737 -38
rect 799 38 833 54
rect 799 -54 833 -38
rect 895 38 929 54
rect 895 -54 929 -38
rect 991 38 1025 54
rect 991 -54 1025 -38
rect 1087 38 1121 54
rect 1087 -54 1121 -38
rect 1183 38 1217 54
rect 1183 -54 1217 -38
rect 1279 38 1313 54
rect 1279 -54 1313 -38
rect -1427 -190 -1393 -128
rect 1393 -190 1427 -128
rect -1427 -224 -1331 -190
rect 1331 -224 1427 -190
<< viali >>
rect -1283 88 -1249 122
rect -1150 88 -1057 122
rect -949 88 -299 122
rect -181 88 1237 122
rect -1313 -38 -1279 38
rect -1217 -38 -1183 38
rect -1121 -38 -1087 38
rect -1025 -38 -991 38
rect -929 -38 -895 38
rect -833 -38 -799 38
rect -737 -38 -703 38
rect -641 -38 -607 38
rect -545 -38 -511 38
rect -449 -38 -415 38
rect -353 -38 -319 38
rect -257 -38 -223 38
rect -161 -38 -127 38
rect -65 -38 -31 38
rect 31 -38 65 38
rect 127 -38 161 38
rect 223 -38 257 38
rect 319 -38 353 38
rect 415 -38 449 38
rect 511 -38 545 38
rect 607 -38 641 38
rect 703 -38 737 38
rect 799 -38 833 38
rect 895 -38 929 38
rect 991 -38 1025 38
rect 1087 -38 1121 38
rect 1183 -38 1217 38
rect 1279 -38 1313 38
<< metal1 >>
rect -1295 122 -1237 128
rect -1295 88 -1283 122
rect -1249 88 -1237 122
rect -1295 82 -1237 88
rect -1167 122 -1041 128
rect -1167 88 -1150 122
rect -1057 88 -1041 122
rect -1167 82 -1041 88
rect -975 122 -273 128
rect -975 88 -949 122
rect -299 88 -273 122
rect -975 82 -273 88
rect -207 122 1263 128
rect -207 88 -181 122
rect 1237 88 1263 122
rect -207 82 1263 88
rect -1319 38 -1273 50
rect -1319 -38 -1313 38
rect -1279 -38 -1273 38
rect -1319 -50 -1273 -38
rect -1223 38 -1177 50
rect -1223 -38 -1217 38
rect -1183 -38 -1177 38
rect -1223 -50 -1177 -38
rect -1127 38 -1081 50
rect -1127 -38 -1121 38
rect -1087 -38 -1081 38
rect -1127 -50 -1081 -38
rect -1031 38 -985 50
rect -1031 -38 -1025 38
rect -991 -38 -985 38
rect -1031 -50 -985 -38
rect -935 38 -889 50
rect -935 -38 -929 38
rect -895 -38 -889 38
rect -935 -50 -889 -38
rect -839 38 -793 50
rect -839 -38 -833 38
rect -799 -38 -793 38
rect -839 -50 -793 -38
rect -743 38 -697 50
rect -743 -38 -737 38
rect -703 -38 -697 38
rect -743 -50 -697 -38
rect -647 38 -601 50
rect -647 -38 -641 38
rect -607 -38 -601 38
rect -647 -50 -601 -38
rect -551 38 -505 50
rect -551 -38 -545 38
rect -511 -38 -505 38
rect -551 -50 -505 -38
rect -455 38 -409 50
rect -455 -38 -449 38
rect -415 -38 -409 38
rect -455 -50 -409 -38
rect -359 38 -313 50
rect -359 -38 -353 38
rect -319 -38 -313 38
rect -359 -50 -313 -38
rect -263 38 -217 50
rect -263 -38 -257 38
rect -223 -38 -217 38
rect -263 -50 -217 -38
rect -167 38 -121 50
rect -167 -38 -161 38
rect -127 -38 -121 38
rect -167 -50 -121 -38
rect -71 38 -25 50
rect -71 -38 -65 38
rect -31 -38 -25 38
rect -71 -50 -25 -38
rect 25 38 71 50
rect 25 -38 31 38
rect 65 -38 71 38
rect 25 -50 71 -38
rect 121 38 167 50
rect 121 -38 127 38
rect 161 -38 167 38
rect 121 -50 167 -38
rect 217 38 263 50
rect 217 -38 223 38
rect 257 -38 263 38
rect 217 -50 263 -38
rect 313 38 359 50
rect 313 -38 319 38
rect 353 -38 359 38
rect 313 -50 359 -38
rect 409 38 455 50
rect 409 -38 415 38
rect 449 -38 455 38
rect 409 -50 455 -38
rect 505 38 551 50
rect 505 -38 511 38
rect 545 -38 551 38
rect 505 -50 551 -38
rect 601 38 647 50
rect 601 -38 607 38
rect 641 -38 647 38
rect 601 -50 647 -38
rect 697 38 743 50
rect 697 -38 703 38
rect 737 -38 743 38
rect 697 -50 743 -38
rect 793 38 839 50
rect 793 -38 799 38
rect 833 -38 839 38
rect 793 -50 839 -38
rect 889 38 935 50
rect 889 -38 895 38
rect 929 -38 935 38
rect 889 -50 935 -38
rect 985 38 1031 50
rect 985 -38 991 38
rect 1025 -38 1031 38
rect 985 -50 1031 -38
rect 1081 38 1127 50
rect 1081 -38 1087 38
rect 1121 -38 1127 38
rect 1081 -50 1127 -38
rect 1177 38 1223 50
rect 1177 -38 1183 38
rect 1217 -38 1223 38
rect 1177 -50 1223 -38
rect 1273 38 1319 50
rect 1273 -38 1279 38
rect 1313 -38 1319 38
rect 1273 -50 1319 -38
<< properties >>
string FIXED_BBOX -1410 -207 1410 207
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.15 m 1 nf 27 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
