magic
tech sky130A
magscale 1 2
timestamp 1717363523
<< error_p >>
rect -29 2507 29 2513
rect -29 2473 -17 2507
rect -29 2467 29 2473
rect -29 2297 29 2303
rect -29 2263 -17 2297
rect -29 2257 29 2263
rect -29 2189 29 2195
rect -29 2155 -17 2189
rect -29 2149 29 2155
rect -29 1979 29 1985
rect -29 1945 -17 1979
rect -29 1939 29 1945
rect -29 1871 29 1877
rect -29 1837 -17 1871
rect -29 1831 29 1837
rect -29 1661 29 1667
rect -29 1627 -17 1661
rect -29 1621 29 1627
rect -29 1553 29 1559
rect -29 1519 -17 1553
rect -29 1513 29 1519
rect -29 1343 29 1349
rect -29 1309 -17 1343
rect -29 1303 29 1309
rect -29 1235 29 1241
rect -29 1201 -17 1235
rect -29 1195 29 1201
rect -29 1025 29 1031
rect -29 991 -17 1025
rect -29 985 29 991
rect -29 917 29 923
rect -29 883 -17 917
rect -29 877 29 883
rect -29 707 29 713
rect -29 673 -17 707
rect -29 667 29 673
rect -29 599 29 605
rect -29 565 -17 599
rect -29 559 29 565
rect -29 389 29 395
rect -29 355 -17 389
rect -29 349 29 355
rect -29 281 29 287
rect -29 247 -17 281
rect -29 241 29 247
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -247 29 -241
rect -29 -281 -17 -247
rect -29 -287 29 -281
rect -29 -355 29 -349
rect -29 -389 -17 -355
rect -29 -395 29 -389
rect -29 -565 29 -559
rect -29 -599 -17 -565
rect -29 -605 29 -599
rect -29 -673 29 -667
rect -29 -707 -17 -673
rect -29 -713 29 -707
rect -29 -883 29 -877
rect -29 -917 -17 -883
rect -29 -923 29 -917
rect -29 -991 29 -985
rect -29 -1025 -17 -991
rect -29 -1031 29 -1025
rect -29 -1201 29 -1195
rect -29 -1235 -17 -1201
rect -29 -1241 29 -1235
rect -29 -1309 29 -1303
rect -29 -1343 -17 -1309
rect -29 -1349 29 -1343
rect -29 -1519 29 -1513
rect -29 -1553 -17 -1519
rect -29 -1559 29 -1553
rect -29 -1627 29 -1621
rect -29 -1661 -17 -1627
rect -29 -1667 29 -1661
rect -29 -1837 29 -1831
rect -29 -1871 -17 -1837
rect -29 -1877 29 -1871
rect -29 -1945 29 -1939
rect -29 -1979 -17 -1945
rect -29 -1985 29 -1979
rect -29 -2155 29 -2149
rect -29 -2189 -17 -2155
rect -29 -2195 29 -2189
rect -29 -2263 29 -2257
rect -29 -2297 -17 -2263
rect -29 -2303 29 -2297
rect -29 -2473 29 -2467
rect -29 -2507 -17 -2473
rect -29 -2513 29 -2507
<< pwell >>
rect -211 -2645 211 2645
<< nmos >>
rect -15 2335 15 2435
rect -15 2017 15 2117
rect -15 1699 15 1799
rect -15 1381 15 1481
rect -15 1063 15 1163
rect -15 745 15 845
rect -15 427 15 527
rect -15 109 15 209
rect -15 -209 15 -109
rect -15 -527 15 -427
rect -15 -845 15 -745
rect -15 -1163 15 -1063
rect -15 -1481 15 -1381
rect -15 -1799 15 -1699
rect -15 -2117 15 -2017
rect -15 -2435 15 -2335
<< ndiff >>
rect -73 2423 -15 2435
rect -73 2347 -61 2423
rect -27 2347 -15 2423
rect -73 2335 -15 2347
rect 15 2423 73 2435
rect 15 2347 27 2423
rect 61 2347 73 2423
rect 15 2335 73 2347
rect -73 2105 -15 2117
rect -73 2029 -61 2105
rect -27 2029 -15 2105
rect -73 2017 -15 2029
rect 15 2105 73 2117
rect 15 2029 27 2105
rect 61 2029 73 2105
rect 15 2017 73 2029
rect -73 1787 -15 1799
rect -73 1711 -61 1787
rect -27 1711 -15 1787
rect -73 1699 -15 1711
rect 15 1787 73 1799
rect 15 1711 27 1787
rect 61 1711 73 1787
rect 15 1699 73 1711
rect -73 1469 -15 1481
rect -73 1393 -61 1469
rect -27 1393 -15 1469
rect -73 1381 -15 1393
rect 15 1469 73 1481
rect 15 1393 27 1469
rect 61 1393 73 1469
rect 15 1381 73 1393
rect -73 1151 -15 1163
rect -73 1075 -61 1151
rect -27 1075 -15 1151
rect -73 1063 -15 1075
rect 15 1151 73 1163
rect 15 1075 27 1151
rect 61 1075 73 1151
rect 15 1063 73 1075
rect -73 833 -15 845
rect -73 757 -61 833
rect -27 757 -15 833
rect -73 745 -15 757
rect 15 833 73 845
rect 15 757 27 833
rect 61 757 73 833
rect 15 745 73 757
rect -73 515 -15 527
rect -73 439 -61 515
rect -27 439 -15 515
rect -73 427 -15 439
rect 15 515 73 527
rect 15 439 27 515
rect 61 439 73 515
rect 15 427 73 439
rect -73 197 -15 209
rect -73 121 -61 197
rect -27 121 -15 197
rect -73 109 -15 121
rect 15 197 73 209
rect 15 121 27 197
rect 61 121 73 197
rect 15 109 73 121
rect -73 -121 -15 -109
rect -73 -197 -61 -121
rect -27 -197 -15 -121
rect -73 -209 -15 -197
rect 15 -121 73 -109
rect 15 -197 27 -121
rect 61 -197 73 -121
rect 15 -209 73 -197
rect -73 -439 -15 -427
rect -73 -515 -61 -439
rect -27 -515 -15 -439
rect -73 -527 -15 -515
rect 15 -439 73 -427
rect 15 -515 27 -439
rect 61 -515 73 -439
rect 15 -527 73 -515
rect -73 -757 -15 -745
rect -73 -833 -61 -757
rect -27 -833 -15 -757
rect -73 -845 -15 -833
rect 15 -757 73 -745
rect 15 -833 27 -757
rect 61 -833 73 -757
rect 15 -845 73 -833
rect -73 -1075 -15 -1063
rect -73 -1151 -61 -1075
rect -27 -1151 -15 -1075
rect -73 -1163 -15 -1151
rect 15 -1075 73 -1063
rect 15 -1151 27 -1075
rect 61 -1151 73 -1075
rect 15 -1163 73 -1151
rect -73 -1393 -15 -1381
rect -73 -1469 -61 -1393
rect -27 -1469 -15 -1393
rect -73 -1481 -15 -1469
rect 15 -1393 73 -1381
rect 15 -1469 27 -1393
rect 61 -1469 73 -1393
rect 15 -1481 73 -1469
rect -73 -1711 -15 -1699
rect -73 -1787 -61 -1711
rect -27 -1787 -15 -1711
rect -73 -1799 -15 -1787
rect 15 -1711 73 -1699
rect 15 -1787 27 -1711
rect 61 -1787 73 -1711
rect 15 -1799 73 -1787
rect -73 -2029 -15 -2017
rect -73 -2105 -61 -2029
rect -27 -2105 -15 -2029
rect -73 -2117 -15 -2105
rect 15 -2029 73 -2017
rect 15 -2105 27 -2029
rect 61 -2105 73 -2029
rect 15 -2117 73 -2105
rect -73 -2347 -15 -2335
rect -73 -2423 -61 -2347
rect -27 -2423 -15 -2347
rect -73 -2435 -15 -2423
rect 15 -2347 73 -2335
rect 15 -2423 27 -2347
rect 61 -2423 73 -2347
rect 15 -2435 73 -2423
<< ndiffc >>
rect -61 2347 -27 2423
rect 27 2347 61 2423
rect -61 2029 -27 2105
rect 27 2029 61 2105
rect -61 1711 -27 1787
rect 27 1711 61 1787
rect -61 1393 -27 1469
rect 27 1393 61 1469
rect -61 1075 -27 1151
rect 27 1075 61 1151
rect -61 757 -27 833
rect 27 757 61 833
rect -61 439 -27 515
rect 27 439 61 515
rect -61 121 -27 197
rect 27 121 61 197
rect -61 -197 -27 -121
rect 27 -197 61 -121
rect -61 -515 -27 -439
rect 27 -515 61 -439
rect -61 -833 -27 -757
rect 27 -833 61 -757
rect -61 -1151 -27 -1075
rect 27 -1151 61 -1075
rect -61 -1469 -27 -1393
rect 27 -1469 61 -1393
rect -61 -1787 -27 -1711
rect 27 -1787 61 -1711
rect -61 -2105 -27 -2029
rect 27 -2105 61 -2029
rect -61 -2423 -27 -2347
rect 27 -2423 61 -2347
<< psubdiff >>
rect -175 2575 -79 2609
rect 79 2575 175 2609
rect -175 2513 -141 2575
rect 141 2513 175 2575
rect -175 -2575 -141 -2513
rect 141 -2575 175 -2513
rect -175 -2609 -79 -2575
rect 79 -2609 175 -2575
<< psubdiffcont >>
rect -79 2575 79 2609
rect -175 -2513 -141 2513
rect 141 -2513 175 2513
rect -79 -2609 79 -2575
<< poly >>
rect -33 2507 33 2523
rect -33 2473 -17 2507
rect 17 2473 33 2507
rect -33 2457 33 2473
rect -15 2435 15 2457
rect -15 2313 15 2335
rect -33 2297 33 2313
rect -33 2263 -17 2297
rect 17 2263 33 2297
rect -33 2247 33 2263
rect -33 2189 33 2205
rect -33 2155 -17 2189
rect 17 2155 33 2189
rect -33 2139 33 2155
rect -15 2117 15 2139
rect -15 1995 15 2017
rect -33 1979 33 1995
rect -33 1945 -17 1979
rect 17 1945 33 1979
rect -33 1929 33 1945
rect -33 1871 33 1887
rect -33 1837 -17 1871
rect 17 1837 33 1871
rect -33 1821 33 1837
rect -15 1799 15 1821
rect -15 1677 15 1699
rect -33 1661 33 1677
rect -33 1627 -17 1661
rect 17 1627 33 1661
rect -33 1611 33 1627
rect -33 1553 33 1569
rect -33 1519 -17 1553
rect 17 1519 33 1553
rect -33 1503 33 1519
rect -15 1481 15 1503
rect -15 1359 15 1381
rect -33 1343 33 1359
rect -33 1309 -17 1343
rect 17 1309 33 1343
rect -33 1293 33 1309
rect -33 1235 33 1251
rect -33 1201 -17 1235
rect 17 1201 33 1235
rect -33 1185 33 1201
rect -15 1163 15 1185
rect -15 1041 15 1063
rect -33 1025 33 1041
rect -33 991 -17 1025
rect 17 991 33 1025
rect -33 975 33 991
rect -33 917 33 933
rect -33 883 -17 917
rect 17 883 33 917
rect -33 867 33 883
rect -15 845 15 867
rect -15 723 15 745
rect -33 707 33 723
rect -33 673 -17 707
rect 17 673 33 707
rect -33 657 33 673
rect -33 599 33 615
rect -33 565 -17 599
rect 17 565 33 599
rect -33 549 33 565
rect -15 527 15 549
rect -15 405 15 427
rect -33 389 33 405
rect -33 355 -17 389
rect 17 355 33 389
rect -33 339 33 355
rect -33 281 33 297
rect -33 247 -17 281
rect 17 247 33 281
rect -33 231 33 247
rect -15 209 15 231
rect -15 87 15 109
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -109 15 -87
rect -15 -231 15 -209
rect -33 -247 33 -231
rect -33 -281 -17 -247
rect 17 -281 33 -247
rect -33 -297 33 -281
rect -33 -355 33 -339
rect -33 -389 -17 -355
rect 17 -389 33 -355
rect -33 -405 33 -389
rect -15 -427 15 -405
rect -15 -549 15 -527
rect -33 -565 33 -549
rect -33 -599 -17 -565
rect 17 -599 33 -565
rect -33 -615 33 -599
rect -33 -673 33 -657
rect -33 -707 -17 -673
rect 17 -707 33 -673
rect -33 -723 33 -707
rect -15 -745 15 -723
rect -15 -867 15 -845
rect -33 -883 33 -867
rect -33 -917 -17 -883
rect 17 -917 33 -883
rect -33 -933 33 -917
rect -33 -991 33 -975
rect -33 -1025 -17 -991
rect 17 -1025 33 -991
rect -33 -1041 33 -1025
rect -15 -1063 15 -1041
rect -15 -1185 15 -1163
rect -33 -1201 33 -1185
rect -33 -1235 -17 -1201
rect 17 -1235 33 -1201
rect -33 -1251 33 -1235
rect -33 -1309 33 -1293
rect -33 -1343 -17 -1309
rect 17 -1343 33 -1309
rect -33 -1359 33 -1343
rect -15 -1381 15 -1359
rect -15 -1503 15 -1481
rect -33 -1519 33 -1503
rect -33 -1553 -17 -1519
rect 17 -1553 33 -1519
rect -33 -1569 33 -1553
rect -33 -1627 33 -1611
rect -33 -1661 -17 -1627
rect 17 -1661 33 -1627
rect -33 -1677 33 -1661
rect -15 -1699 15 -1677
rect -15 -1821 15 -1799
rect -33 -1837 33 -1821
rect -33 -1871 -17 -1837
rect 17 -1871 33 -1837
rect -33 -1887 33 -1871
rect -33 -1945 33 -1929
rect -33 -1979 -17 -1945
rect 17 -1979 33 -1945
rect -33 -1995 33 -1979
rect -15 -2017 15 -1995
rect -15 -2139 15 -2117
rect -33 -2155 33 -2139
rect -33 -2189 -17 -2155
rect 17 -2189 33 -2155
rect -33 -2205 33 -2189
rect -33 -2263 33 -2247
rect -33 -2297 -17 -2263
rect 17 -2297 33 -2263
rect -33 -2313 33 -2297
rect -15 -2335 15 -2313
rect -15 -2457 15 -2435
rect -33 -2473 33 -2457
rect -33 -2507 -17 -2473
rect 17 -2507 33 -2473
rect -33 -2523 33 -2507
<< polycont >>
rect -17 2473 17 2507
rect -17 2263 17 2297
rect -17 2155 17 2189
rect -17 1945 17 1979
rect -17 1837 17 1871
rect -17 1627 17 1661
rect -17 1519 17 1553
rect -17 1309 17 1343
rect -17 1201 17 1235
rect -17 991 17 1025
rect -17 883 17 917
rect -17 673 17 707
rect -17 565 17 599
rect -17 355 17 389
rect -17 247 17 281
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -281 17 -247
rect -17 -389 17 -355
rect -17 -599 17 -565
rect -17 -707 17 -673
rect -17 -917 17 -883
rect -17 -1025 17 -991
rect -17 -1235 17 -1201
rect -17 -1343 17 -1309
rect -17 -1553 17 -1519
rect -17 -1661 17 -1627
rect -17 -1871 17 -1837
rect -17 -1979 17 -1945
rect -17 -2189 17 -2155
rect -17 -2297 17 -2263
rect -17 -2507 17 -2473
<< locali >>
rect -175 2575 -79 2609
rect 79 2575 175 2609
rect -175 2513 -141 2575
rect 141 2513 175 2575
rect -33 2473 -17 2507
rect 17 2473 33 2507
rect -61 2423 -27 2439
rect -61 2331 -27 2347
rect 27 2423 61 2439
rect 27 2331 61 2347
rect -33 2263 -17 2297
rect 17 2263 33 2297
rect -33 2155 -17 2189
rect 17 2155 33 2189
rect -61 2105 -27 2121
rect -61 2013 -27 2029
rect 27 2105 61 2121
rect 27 2013 61 2029
rect -33 1945 -17 1979
rect 17 1945 33 1979
rect -33 1837 -17 1871
rect 17 1837 33 1871
rect -61 1787 -27 1803
rect -61 1695 -27 1711
rect 27 1787 61 1803
rect 27 1695 61 1711
rect -33 1627 -17 1661
rect 17 1627 33 1661
rect -33 1519 -17 1553
rect 17 1519 33 1553
rect -61 1469 -27 1485
rect -61 1377 -27 1393
rect 27 1469 61 1485
rect 27 1377 61 1393
rect -33 1309 -17 1343
rect 17 1309 33 1343
rect -33 1201 -17 1235
rect 17 1201 33 1235
rect -61 1151 -27 1167
rect -61 1059 -27 1075
rect 27 1151 61 1167
rect 27 1059 61 1075
rect -33 991 -17 1025
rect 17 991 33 1025
rect -33 883 -17 917
rect 17 883 33 917
rect -61 833 -27 849
rect -61 741 -27 757
rect 27 833 61 849
rect 27 741 61 757
rect -33 673 -17 707
rect 17 673 33 707
rect -33 565 -17 599
rect 17 565 33 599
rect -61 515 -27 531
rect -61 423 -27 439
rect 27 515 61 531
rect 27 423 61 439
rect -33 355 -17 389
rect 17 355 33 389
rect -33 247 -17 281
rect 17 247 33 281
rect -61 197 -27 213
rect -61 105 -27 121
rect 27 197 61 213
rect 27 105 61 121
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -121 -27 -105
rect -61 -213 -27 -197
rect 27 -121 61 -105
rect 27 -213 61 -197
rect -33 -281 -17 -247
rect 17 -281 33 -247
rect -33 -389 -17 -355
rect 17 -389 33 -355
rect -61 -439 -27 -423
rect -61 -531 -27 -515
rect 27 -439 61 -423
rect 27 -531 61 -515
rect -33 -599 -17 -565
rect 17 -599 33 -565
rect -33 -707 -17 -673
rect 17 -707 33 -673
rect -61 -757 -27 -741
rect -61 -849 -27 -833
rect 27 -757 61 -741
rect 27 -849 61 -833
rect -33 -917 -17 -883
rect 17 -917 33 -883
rect -33 -1025 -17 -991
rect 17 -1025 33 -991
rect -61 -1075 -27 -1059
rect -61 -1167 -27 -1151
rect 27 -1075 61 -1059
rect 27 -1167 61 -1151
rect -33 -1235 -17 -1201
rect 17 -1235 33 -1201
rect -33 -1343 -17 -1309
rect 17 -1343 33 -1309
rect -61 -1393 -27 -1377
rect -61 -1485 -27 -1469
rect 27 -1393 61 -1377
rect 27 -1485 61 -1469
rect -33 -1553 -17 -1519
rect 17 -1553 33 -1519
rect -33 -1661 -17 -1627
rect 17 -1661 33 -1627
rect -61 -1711 -27 -1695
rect -61 -1803 -27 -1787
rect 27 -1711 61 -1695
rect 27 -1803 61 -1787
rect -33 -1871 -17 -1837
rect 17 -1871 33 -1837
rect -33 -1979 -17 -1945
rect 17 -1979 33 -1945
rect -61 -2029 -27 -2013
rect -61 -2121 -27 -2105
rect 27 -2029 61 -2013
rect 27 -2121 61 -2105
rect -33 -2189 -17 -2155
rect 17 -2189 33 -2155
rect -33 -2297 -17 -2263
rect 17 -2297 33 -2263
rect -61 -2347 -27 -2331
rect -61 -2439 -27 -2423
rect 27 -2347 61 -2331
rect 27 -2439 61 -2423
rect -33 -2507 -17 -2473
rect 17 -2507 33 -2473
rect -175 -2575 -141 -2513
rect 141 -2575 175 -2513
rect -175 -2609 -79 -2575
rect 79 -2609 175 -2575
<< viali >>
rect -17 2473 17 2507
rect -61 2347 -27 2423
rect 27 2347 61 2423
rect -17 2263 17 2297
rect -17 2155 17 2189
rect -61 2029 -27 2105
rect 27 2029 61 2105
rect -17 1945 17 1979
rect -17 1837 17 1871
rect -61 1711 -27 1787
rect 27 1711 61 1787
rect -17 1627 17 1661
rect -17 1519 17 1553
rect -61 1393 -27 1469
rect 27 1393 61 1469
rect -17 1309 17 1343
rect -17 1201 17 1235
rect -61 1075 -27 1151
rect 27 1075 61 1151
rect -17 991 17 1025
rect -17 883 17 917
rect -61 757 -27 833
rect 27 757 61 833
rect -17 673 17 707
rect -17 565 17 599
rect -61 439 -27 515
rect 27 439 61 515
rect -17 355 17 389
rect -17 247 17 281
rect -61 121 -27 197
rect 27 121 61 197
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -197 -27 -121
rect 27 -197 61 -121
rect -17 -281 17 -247
rect -17 -389 17 -355
rect -61 -515 -27 -439
rect 27 -515 61 -439
rect -17 -599 17 -565
rect -17 -707 17 -673
rect -61 -833 -27 -757
rect 27 -833 61 -757
rect -17 -917 17 -883
rect -17 -1025 17 -991
rect -61 -1151 -27 -1075
rect 27 -1151 61 -1075
rect -17 -1235 17 -1201
rect -17 -1343 17 -1309
rect -61 -1469 -27 -1393
rect 27 -1469 61 -1393
rect -17 -1553 17 -1519
rect -17 -1661 17 -1627
rect -61 -1787 -27 -1711
rect 27 -1787 61 -1711
rect -17 -1871 17 -1837
rect -17 -1979 17 -1945
rect -61 -2105 -27 -2029
rect 27 -2105 61 -2029
rect -17 -2189 17 -2155
rect -17 -2297 17 -2263
rect -61 -2423 -27 -2347
rect 27 -2423 61 -2347
rect -17 -2507 17 -2473
<< metal1 >>
rect -29 2507 29 2513
rect -29 2473 -17 2507
rect 17 2473 29 2507
rect -29 2467 29 2473
rect -67 2423 -21 2435
rect -67 2347 -61 2423
rect -27 2347 -21 2423
rect -67 2335 -21 2347
rect 21 2423 67 2435
rect 21 2347 27 2423
rect 61 2347 67 2423
rect 21 2335 67 2347
rect -29 2297 29 2303
rect -29 2263 -17 2297
rect 17 2263 29 2297
rect -29 2257 29 2263
rect -29 2189 29 2195
rect -29 2155 -17 2189
rect 17 2155 29 2189
rect -29 2149 29 2155
rect -67 2105 -21 2117
rect -67 2029 -61 2105
rect -27 2029 -21 2105
rect -67 2017 -21 2029
rect 21 2105 67 2117
rect 21 2029 27 2105
rect 61 2029 67 2105
rect 21 2017 67 2029
rect -29 1979 29 1985
rect -29 1945 -17 1979
rect 17 1945 29 1979
rect -29 1939 29 1945
rect -29 1871 29 1877
rect -29 1837 -17 1871
rect 17 1837 29 1871
rect -29 1831 29 1837
rect -67 1787 -21 1799
rect -67 1711 -61 1787
rect -27 1711 -21 1787
rect -67 1699 -21 1711
rect 21 1787 67 1799
rect 21 1711 27 1787
rect 61 1711 67 1787
rect 21 1699 67 1711
rect -29 1661 29 1667
rect -29 1627 -17 1661
rect 17 1627 29 1661
rect -29 1621 29 1627
rect -29 1553 29 1559
rect -29 1519 -17 1553
rect 17 1519 29 1553
rect -29 1513 29 1519
rect -67 1469 -21 1481
rect -67 1393 -61 1469
rect -27 1393 -21 1469
rect -67 1381 -21 1393
rect 21 1469 67 1481
rect 21 1393 27 1469
rect 61 1393 67 1469
rect 21 1381 67 1393
rect -29 1343 29 1349
rect -29 1309 -17 1343
rect 17 1309 29 1343
rect -29 1303 29 1309
rect -29 1235 29 1241
rect -29 1201 -17 1235
rect 17 1201 29 1235
rect -29 1195 29 1201
rect -67 1151 -21 1163
rect -67 1075 -61 1151
rect -27 1075 -21 1151
rect -67 1063 -21 1075
rect 21 1151 67 1163
rect 21 1075 27 1151
rect 61 1075 67 1151
rect 21 1063 67 1075
rect -29 1025 29 1031
rect -29 991 -17 1025
rect 17 991 29 1025
rect -29 985 29 991
rect -29 917 29 923
rect -29 883 -17 917
rect 17 883 29 917
rect -29 877 29 883
rect -67 833 -21 845
rect -67 757 -61 833
rect -27 757 -21 833
rect -67 745 -21 757
rect 21 833 67 845
rect 21 757 27 833
rect 61 757 67 833
rect 21 745 67 757
rect -29 707 29 713
rect -29 673 -17 707
rect 17 673 29 707
rect -29 667 29 673
rect -29 599 29 605
rect -29 565 -17 599
rect 17 565 29 599
rect -29 559 29 565
rect -67 515 -21 527
rect -67 439 -61 515
rect -27 439 -21 515
rect -67 427 -21 439
rect 21 515 67 527
rect 21 439 27 515
rect 61 439 67 515
rect 21 427 67 439
rect -29 389 29 395
rect -29 355 -17 389
rect 17 355 29 389
rect -29 349 29 355
rect -29 281 29 287
rect -29 247 -17 281
rect 17 247 29 281
rect -29 241 29 247
rect -67 197 -21 209
rect -67 121 -61 197
rect -27 121 -21 197
rect -67 109 -21 121
rect 21 197 67 209
rect 21 121 27 197
rect 61 121 67 197
rect 21 109 67 121
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -121 -21 -109
rect -67 -197 -61 -121
rect -27 -197 -21 -121
rect -67 -209 -21 -197
rect 21 -121 67 -109
rect 21 -197 27 -121
rect 61 -197 67 -121
rect 21 -209 67 -197
rect -29 -247 29 -241
rect -29 -281 -17 -247
rect 17 -281 29 -247
rect -29 -287 29 -281
rect -29 -355 29 -349
rect -29 -389 -17 -355
rect 17 -389 29 -355
rect -29 -395 29 -389
rect -67 -439 -21 -427
rect -67 -515 -61 -439
rect -27 -515 -21 -439
rect -67 -527 -21 -515
rect 21 -439 67 -427
rect 21 -515 27 -439
rect 61 -515 67 -439
rect 21 -527 67 -515
rect -29 -565 29 -559
rect -29 -599 -17 -565
rect 17 -599 29 -565
rect -29 -605 29 -599
rect -29 -673 29 -667
rect -29 -707 -17 -673
rect 17 -707 29 -673
rect -29 -713 29 -707
rect -67 -757 -21 -745
rect -67 -833 -61 -757
rect -27 -833 -21 -757
rect -67 -845 -21 -833
rect 21 -757 67 -745
rect 21 -833 27 -757
rect 61 -833 67 -757
rect 21 -845 67 -833
rect -29 -883 29 -877
rect -29 -917 -17 -883
rect 17 -917 29 -883
rect -29 -923 29 -917
rect -29 -991 29 -985
rect -29 -1025 -17 -991
rect 17 -1025 29 -991
rect -29 -1031 29 -1025
rect -67 -1075 -21 -1063
rect -67 -1151 -61 -1075
rect -27 -1151 -21 -1075
rect -67 -1163 -21 -1151
rect 21 -1075 67 -1063
rect 21 -1151 27 -1075
rect 61 -1151 67 -1075
rect 21 -1163 67 -1151
rect -29 -1201 29 -1195
rect -29 -1235 -17 -1201
rect 17 -1235 29 -1201
rect -29 -1241 29 -1235
rect -29 -1309 29 -1303
rect -29 -1343 -17 -1309
rect 17 -1343 29 -1309
rect -29 -1349 29 -1343
rect -67 -1393 -21 -1381
rect -67 -1469 -61 -1393
rect -27 -1469 -21 -1393
rect -67 -1481 -21 -1469
rect 21 -1393 67 -1381
rect 21 -1469 27 -1393
rect 61 -1469 67 -1393
rect 21 -1481 67 -1469
rect -29 -1519 29 -1513
rect -29 -1553 -17 -1519
rect 17 -1553 29 -1519
rect -29 -1559 29 -1553
rect -29 -1627 29 -1621
rect -29 -1661 -17 -1627
rect 17 -1661 29 -1627
rect -29 -1667 29 -1661
rect -67 -1711 -21 -1699
rect -67 -1787 -61 -1711
rect -27 -1787 -21 -1711
rect -67 -1799 -21 -1787
rect 21 -1711 67 -1699
rect 21 -1787 27 -1711
rect 61 -1787 67 -1711
rect 21 -1799 67 -1787
rect -29 -1837 29 -1831
rect -29 -1871 -17 -1837
rect 17 -1871 29 -1837
rect -29 -1877 29 -1871
rect -29 -1945 29 -1939
rect -29 -1979 -17 -1945
rect 17 -1979 29 -1945
rect -29 -1985 29 -1979
rect -67 -2029 -21 -2017
rect -67 -2105 -61 -2029
rect -27 -2105 -21 -2029
rect -67 -2117 -21 -2105
rect 21 -2029 67 -2017
rect 21 -2105 27 -2029
rect 61 -2105 67 -2029
rect 21 -2117 67 -2105
rect -29 -2155 29 -2149
rect -29 -2189 -17 -2155
rect 17 -2189 29 -2155
rect -29 -2195 29 -2189
rect -29 -2263 29 -2257
rect -29 -2297 -17 -2263
rect 17 -2297 29 -2263
rect -29 -2303 29 -2297
rect -67 -2347 -21 -2335
rect -67 -2423 -61 -2347
rect -27 -2423 -21 -2347
rect -67 -2435 -21 -2423
rect 21 -2347 67 -2335
rect 21 -2423 27 -2347
rect 61 -2423 67 -2347
rect 21 -2435 67 -2423
rect -29 -2473 29 -2467
rect -29 -2507 -17 -2473
rect 17 -2507 29 -2473
rect -29 -2513 29 -2507
<< properties >>
string FIXED_BBOX -158 -2592 158 2592
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.15 m 16 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
