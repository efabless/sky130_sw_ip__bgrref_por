magic
tech sky130A
magscale 1 2
timestamp 1717527227
<< nwell >>
rect -263 -477 263 477
<< pmos >>
rect -63 118 -33 258
rect 33 118 63 258
rect -63 -258 -33 -118
rect 33 -258 63 -118
<< pdiff >>
rect -125 246 -63 258
rect -125 130 -113 246
rect -79 130 -63 246
rect -125 118 -63 130
rect -33 246 33 258
rect -33 130 -17 246
rect 17 130 33 246
rect -33 118 33 130
rect 63 246 125 258
rect 63 130 79 246
rect 113 130 125 246
rect 63 118 125 130
rect -125 -130 -63 -118
rect -125 -246 -113 -130
rect -79 -246 -63 -130
rect -125 -258 -63 -246
rect -33 -130 33 -118
rect -33 -246 -17 -130
rect 17 -246 33 -130
rect -33 -258 33 -246
rect 63 -130 125 -118
rect 63 -246 79 -130
rect 113 -246 125 -130
rect 63 -258 125 -246
<< pdiffc >>
rect -113 130 -79 246
rect -17 130 17 246
rect 79 130 113 246
rect -113 -246 -79 -130
rect -17 -246 17 -130
rect 79 -246 113 -130
<< nsubdiff >>
rect -227 407 -131 441
rect 131 407 227 441
rect -227 345 -193 407
rect 193 345 227 407
rect -227 -407 -193 -345
rect 193 -407 227 -345
rect -227 -441 -131 -407
rect 131 -441 227 -407
<< nsubdiffcont >>
rect -131 407 131 441
rect -227 -345 -193 345
rect 193 -345 227 345
rect -131 -441 131 -407
<< poly >>
rect -81 339 81 355
rect -81 305 -65 339
rect -31 305 31 339
rect 65 305 81 339
rect -81 289 81 305
rect -63 258 -33 289
rect 33 258 63 289
rect -63 87 -33 118
rect 33 87 63 118
rect -81 71 81 87
rect -81 37 -65 71
rect -31 37 31 71
rect 65 37 81 71
rect -81 21 81 37
rect -81 -37 81 -21
rect -81 -71 -65 -37
rect -31 -71 31 -37
rect 65 -71 81 -37
rect -81 -87 81 -71
rect -63 -118 -33 -87
rect 33 -118 63 -87
rect -63 -289 -33 -258
rect 33 -289 63 -258
rect -81 -305 81 -289
rect -81 -339 -65 -305
rect -31 -339 31 -305
rect 65 -339 81 -305
rect -81 -355 81 -339
<< polycont >>
rect -65 305 -31 339
rect 31 305 65 339
rect -65 37 -31 71
rect 31 37 65 71
rect -65 -71 -31 -37
rect 31 -71 65 -37
rect -65 -339 -31 -305
rect 31 -339 65 -305
<< locali >>
rect -227 407 -131 441
rect 131 407 227 441
rect -227 345 -193 407
rect 193 345 227 407
rect -81 305 -65 339
rect -31 305 31 339
rect 65 305 81 339
rect -113 246 -79 262
rect -113 114 -79 130
rect -17 246 17 262
rect -17 114 17 130
rect 79 246 113 262
rect 79 114 113 130
rect -81 37 -65 71
rect -31 37 31 71
rect 65 37 81 71
rect -81 -71 -65 -37
rect -31 -71 31 -37
rect 65 -71 81 -37
rect -113 -130 -79 -114
rect -113 -262 -79 -246
rect -17 -130 17 -114
rect -17 -262 17 -246
rect 79 -130 113 -114
rect 79 -262 113 -246
rect -81 -339 -65 -305
rect -31 -339 31 -305
rect 65 -339 81 -305
rect -227 -407 -193 -345
rect 193 -407 227 -345
rect -227 -441 -131 -407
rect 131 -441 227 -407
<< viali >>
rect -65 305 -31 339
rect 31 305 65 339
rect -113 130 -79 246
rect -17 130 17 246
rect 79 130 113 246
rect -65 37 -31 71
rect 31 37 65 71
rect -65 -71 -31 -37
rect 31 -71 65 -37
rect -113 -246 -79 -130
rect -17 -246 17 -130
rect 79 -246 113 -130
rect -65 -339 -31 -305
rect 31 -339 65 -305
<< metal1 >>
rect -77 339 77 345
rect -77 305 -65 339
rect -31 305 31 339
rect 65 305 77 339
rect -77 299 77 305
rect -119 246 -73 258
rect -119 130 -113 246
rect -79 130 -73 246
rect -119 118 -73 130
rect -23 246 23 258
rect -23 130 -17 246
rect 17 130 23 246
rect -23 118 23 130
rect 73 246 119 258
rect 73 130 79 246
rect 113 130 119 246
rect 73 118 119 130
rect -77 71 77 77
rect -77 37 -65 71
rect -31 37 31 71
rect 65 37 77 71
rect -77 31 77 37
rect -77 -37 77 -31
rect -77 -71 -65 -37
rect -31 -71 31 -37
rect 65 -71 77 -37
rect -77 -77 77 -71
rect -119 -130 -73 -118
rect -119 -246 -113 -130
rect -79 -246 -73 -130
rect -119 -258 -73 -246
rect -23 -130 23 -118
rect -23 -246 -17 -130
rect 17 -246 23 -130
rect -23 -258 23 -246
rect 73 -130 119 -118
rect 73 -246 79 -130
rect 113 -246 119 -130
rect 73 -258 119 -246
rect -77 -305 77 -299
rect -77 -339 -65 -305
rect -31 -339 31 -305
rect 65 -339 77 -305
rect -77 -345 77 -339
<< properties >>
string FIXED_BBOX -210 -424 210 424
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.7 l 0.15 m 2 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
