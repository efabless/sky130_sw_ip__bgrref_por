magic
tech sky130A
magscale 1 2
timestamp 1721073345
<< isosubstrate >>
rect 3992 -292617 17571 -285669
<< nwell >>
rect 3668 -285550 38526 -285370
rect 3668 -292646 3908 -285550
rect 38286 -292646 38526 -285550
rect 3668 -292890 38526 -292646
<< mvpsubdiff >>
rect 3489 -285237 3549 -285203
rect 38627 -285237 38687 -285203
rect 3489 -285263 3523 -285237
rect 38653 -285263 38687 -285237
rect 3489 -293013 3523 -292987
rect 38653 -293013 38687 -292987
rect 3489 -293047 3549 -293013
rect 38627 -293047 38687 -293013
<< mvnsubdiff >>
rect 3734 -285470 3794 -285436
rect 38400 -285470 38460 -285436
rect 3734 -285496 3768 -285470
rect 3734 -292790 3768 -292764
rect 38426 -285496 38460 -285470
rect 38426 -292790 38460 -292764
rect 3734 -292824 3794 -292790
rect 38400 -292824 38460 -292790
<< mvpsubdiffcont >>
rect 3549 -285237 38627 -285203
rect 3489 -292987 3523 -285263
rect 38653 -292987 38687 -285263
rect 3549 -293047 38627 -293013
<< mvnsubdiffcont >>
rect 3794 -285470 38400 -285436
rect 3734 -292764 3768 -285496
rect 38426 -292764 38460 -285496
rect 3794 -292824 38400 -292790
<< locali >>
rect 3489 -285237 3549 -285203
rect 38627 -285237 38687 -285203
rect 3489 -285263 38687 -285237
rect 3523 -285274 38653 -285263
rect 3523 -285320 3551 -285274
rect 38510 -285306 38653 -285274
rect 38510 -285320 38595 -285306
rect 3523 -285370 38595 -285320
rect 3523 -285407 3633 -285370
rect 3523 -292843 3540 -285407
rect 3583 -292843 3633 -285407
rect 3734 -285470 3794 -285436
rect 38400 -285470 38460 -285436
rect 3734 -285496 38460 -285470
rect 3768 -285506 38426 -285496
rect 3768 -285550 3804 -285506
rect 38319 -285525 38426 -285506
rect 38319 -285550 38363 -285525
rect 3768 -285590 38363 -285550
rect 3768 -285608 3895 -285590
rect 3768 -292656 3802 -285608
rect 3844 -292656 3895 -285608
rect 7353 -285717 15350 -285714
rect 7292 -285760 15350 -285717
rect 7292 -285801 7498 -285760
rect 7292 -289021 7360 -285801
rect 7412 -285816 7498 -285801
rect 15275 -285816 15350 -285760
rect 7412 -285903 15350 -285816
rect 7412 -288909 7481 -285903
rect 11766 -286000 12544 -285903
rect 11766 -288849 12025 -286000
rect 12322 -288849 12544 -286000
rect 11766 -288909 12544 -288849
rect 15161 -285905 15350 -285903
rect 15161 -288182 15216 -285905
rect 15268 -287795 15350 -285905
rect 15928 -287795 16036 -287790
rect 15268 -287903 16036 -287795
rect 15268 -288182 15414 -287903
rect 15161 -288909 15414 -288182
rect 15928 -288909 16036 -287903
rect 7412 -288987 16036 -288909
rect 7412 -289021 7479 -288987
rect 7292 -289047 7479 -289021
rect 9970 -289013 16036 -288987
rect 9970 -289047 13305 -289013
rect 7292 -289062 13305 -289047
rect 15607 -289062 16036 -289013
rect 7292 -289065 16036 -289062
rect 7292 -289098 11061 -289065
rect 11030 -289118 11061 -289098
rect 13220 -289098 16036 -289065
rect 13220 -289118 13244 -289098
rect 11030 -289355 13244 -289118
rect 3768 -292692 3895 -292656
rect 38324 -292692 38363 -285590
rect 3768 -292732 38363 -292692
rect 3768 -292764 3821 -292732
rect 3734 -292769 3821 -292764
rect 38284 -292746 38363 -292732
rect 38402 -292746 38426 -285525
rect 38284 -292764 38426 -292746
rect 38284 -292769 38460 -292764
rect 3734 -292790 38460 -292769
rect 3734 -292824 3794 -292790
rect 38400 -292824 38460 -292790
rect 3523 -292877 3633 -292843
rect 38553 -292873 38595 -285370
rect 38634 -292873 38653 -285306
rect 38553 -292877 38653 -292873
rect 3523 -292942 38653 -292877
rect 3523 -292981 3593 -292942
rect 38616 -292981 38653 -292942
rect 3523 -292987 38653 -292981
rect 3489 -293013 38687 -292987
rect 3489 -293047 3549 -293013
rect 38627 -293047 38687 -293013
<< viali >>
rect 3551 -285320 38510 -285274
rect 3540 -292843 3583 -285407
rect 3804 -285550 38319 -285506
rect 3802 -292656 3844 -285608
rect 7360 -289021 7412 -285801
rect 7498 -285816 15275 -285760
rect 15216 -288182 15268 -285905
rect 7479 -289047 9970 -288987
rect 13305 -289062 15607 -289013
rect 11061 -289118 13220 -289065
rect 3821 -292769 38284 -292732
rect 38363 -292746 38402 -285525
rect 38595 -292873 38634 -285306
rect 3593 -292981 38616 -292942
<< metal1 >>
rect 3493 -285274 38674 -285210
rect 3493 -285320 3551 -285274
rect 38510 -285306 38674 -285274
rect 38510 -285320 38595 -285306
rect 3493 -285362 38595 -285320
rect 3502 -285407 3612 -285362
rect 3502 -292843 3540 -285407
rect 3583 -292843 3612 -285407
rect 3756 -285457 38440 -285453
rect 3756 -285496 38447 -285457
rect 3756 -285506 16368 -285496
rect 24480 -285506 38447 -285496
rect 3756 -285550 3804 -285506
rect 38319 -285525 38447 -285506
rect 38319 -285550 38363 -285525
rect 3756 -285568 16368 -285550
rect 24480 -285568 38363 -285550
rect 3756 -285579 38363 -285568
rect 3756 -285608 3877 -285579
rect 3756 -289178 3802 -285608
rect 3844 -289178 3877 -285608
rect 7295 -285715 7513 -285713
rect 7295 -285760 15350 -285715
rect 7295 -285801 7498 -285760
rect 7295 -289021 7360 -285801
rect 7412 -285816 7498 -285801
rect 15275 -285816 15350 -285760
rect 7412 -285894 15350 -285816
rect 7412 -285997 7513 -285894
rect 15145 -285905 15350 -285894
rect 7412 -286429 7676 -285997
rect 7772 -286429 8008 -285997
rect 8104 -286429 8340 -285997
rect 8436 -286429 8672 -285997
rect 8768 -286429 9004 -285997
rect 9100 -286429 9336 -285997
rect 9432 -286429 9668 -285997
rect 9764 -286429 10000 -285997
rect 10096 -286429 10332 -285997
rect 10428 -286429 10664 -285997
rect 10760 -286429 10996 -285997
rect 11092 -286429 11328 -285997
rect 11424 -286429 11660 -285997
rect 12125 -286429 12716 -286115
rect 12800 -286429 13038 -285996
rect 13134 -286429 13372 -285996
rect 13468 -286429 13706 -285996
rect 13802 -286429 14040 -285996
rect 14136 -286429 14374 -285996
rect 14470 -286429 14708 -285996
rect 14804 -286429 15042 -285996
rect 7412 -288907 7513 -286429
rect 7606 -288829 7842 -288397
rect 7938 -288829 8174 -288397
rect 8270 -288829 8506 -288397
rect 8602 -288829 8838 -288397
rect 8934 -288829 9170 -288397
rect 9266 -288829 9502 -288397
rect 9598 -288829 9834 -288397
rect 9930 -288829 10166 -288397
rect 10262 -288829 10498 -288397
rect 10594 -288829 10830 -288397
rect 10926 -288829 11162 -288397
rect 11258 -288829 11494 -288397
rect 11588 -288747 12197 -288397
rect 11827 -288868 11874 -288747
rect 7412 -288976 10050 -288907
rect 7412 -289021 7467 -288976
rect 7295 -289052 7467 -289021
rect 10015 -289052 10050 -288976
rect 7295 -289094 10050 -289052
rect 10468 -288915 11874 -288868
rect 7901 -289096 8874 -289094
rect 3756 -289467 3772 -289178
rect 3870 -289467 3877 -289178
rect 10468 -289262 10515 -288915
rect 12407 -288953 12455 -286429
rect 15145 -288182 15216 -285905
rect 15268 -288182 15350 -285905
rect 15145 -288235 15350 -288182
rect 15477 -288394 15543 -288023
rect 15791 -288025 15858 -288023
rect 15579 -288067 15858 -288025
rect 15791 -288340 15858 -288067
rect 15579 -288382 15858 -288340
rect 12634 -288829 12872 -288396
rect 12968 -288829 13206 -288396
rect 13302 -288829 13540 -288396
rect 13636 -288829 13874 -288396
rect 13970 -288829 14208 -288396
rect 14304 -288829 14542 -288396
rect 14638 -288829 14876 -288396
rect 14983 -288829 15543 -288394
rect 15791 -288448 15858 -288382
rect 15579 -288490 15858 -288448
rect 15791 -288762 15858 -288490
rect 15579 -288829 15858 -288762
rect 10784 -289001 12455 -288953
rect 13056 -288976 15663 -288972
rect 10784 -289210 10832 -289001
rect 13056 -289013 13403 -288976
rect 15496 -289013 15663 -288976
rect 13056 -289043 13305 -289013
rect 11027 -289062 13305 -289043
rect 15607 -289062 15663 -289013
rect 11027 -289065 15663 -289062
rect 11027 -289118 11061 -289065
rect 13220 -289092 15663 -289065
rect 13220 -289118 13240 -289092
rect 11027 -289355 13240 -289118
rect 15791 -289266 15858 -288829
rect 3756 -292656 3802 -289467
rect 3844 -292656 3877 -289467
rect 17538 -290701 17586 -289045
rect 16990 -290749 17586 -290701
rect 3986 -292610 17746 -292563
rect 3986 -292611 23772 -292610
rect 3756 -292703 3877 -292656
rect 38334 -292703 38363 -285579
rect 3756 -292732 38363 -292703
rect 3756 -292769 3821 -292732
rect 38284 -292746 38363 -292732
rect 38402 -292746 38447 -285525
rect 38284 -292769 38447 -292746
rect 3756 -292802 38447 -292769
rect 3756 -292805 38380 -292802
rect 3758 -292809 38380 -292805
rect 3502 -292902 3612 -292843
rect 38562 -292873 38595 -285362
rect 38634 -285362 38674 -285306
rect 38634 -292873 38672 -285362
rect 38562 -292902 38672 -292873
rect 3502 -292927 38672 -292902
rect 3502 -292942 17403 -292927
rect 24818 -292942 38672 -292927
rect 3502 -292981 3593 -292942
rect 38616 -292981 38672 -292942
rect 3502 -293001 17403 -292981
rect 24818 -293001 38672 -292981
rect 3502 -293032 38672 -293001
rect 38562 -293043 38672 -293032
<< via1 >>
rect 16368 -285506 24480 -285496
rect 16368 -285550 24480 -285506
rect 16368 -285568 24480 -285550
rect 7467 -288987 10015 -288976
rect 7467 -289047 7479 -288987
rect 7479 -289047 9970 -288987
rect 9970 -289047 10015 -288987
rect 7467 -289052 10015 -289047
rect 3772 -289467 3802 -289178
rect 3802 -289467 3844 -289178
rect 3844 -289467 3870 -289178
rect 13403 -289013 15496 -288976
rect 13403 -289041 15496 -289013
rect 16786 -289428 17380 -289293
rect 5791 -292476 9241 -292342
rect 12676 -292483 16558 -292395
rect 17403 -292942 24818 -292927
rect 17403 -292981 24818 -292942
rect 17403 -293001 24818 -292981
<< metal2 >>
rect 16314 -285496 24531 -285457
rect 16314 -285557 16368 -285496
rect 16312 -285568 16368 -285557
rect 24480 -285568 24531 -285496
rect 16312 -285850 24531 -285568
rect 15937 -288806 16181 -287878
rect 7258 -288976 16181 -288806
rect 7258 -289052 7467 -288976
rect 10015 -289041 13403 -288976
rect 15496 -289041 16181 -288976
rect 10015 -289052 16181 -289041
rect 7258 -289070 16181 -289052
rect 7258 -289072 16078 -289070
rect 3464 -289178 4428 -289169
rect 3464 -289467 3772 -289178
rect 3870 -289467 4428 -289178
rect 3464 -289479 4428 -289467
rect 16312 -289476 16605 -285850
rect 24238 -286408 24531 -285850
rect 39385 -287174 39585 -287137
rect 38048 -287293 39585 -287174
rect 39385 -287337 39585 -287293
rect 16747 -288187 17828 -287923
rect 16747 -289293 17438 -288187
rect 39296 -289256 39496 -289188
rect 16747 -289428 16786 -289293
rect 17380 -289428 17438 -289293
rect 38044 -289340 39496 -289256
rect 39296 -289388 39496 -289340
rect 16747 -289466 17438 -289428
rect 35038 -290006 39195 -290005
rect 35038 -290381 39497 -290006
rect 39301 -290786 39501 -290729
rect 37952 -290871 39501 -290786
rect 37952 -291076 38037 -290871
rect 39301 -290929 39501 -290871
rect 4462 -292342 9298 -292313
rect 3569 -292649 4341 -292449
rect 4462 -292476 5791 -292342
rect 9241 -292476 9298 -292342
rect 4462 -292805 9298 -292476
rect 12630 -292395 16597 -292360
rect 12630 -292483 12676 -292395
rect 16558 -292483 16597 -292395
rect 12630 -292805 16597 -292483
rect 4462 -292806 16600 -292805
rect 3564 -293345 16600 -292806
rect 4462 -293347 16600 -293345
rect 17324 -292927 17872 -292805
rect 17324 -293001 17403 -292927
rect 17324 -293003 17872 -293001
rect 17324 -293338 24877 -293003
rect 17324 -293347 17872 -293338
use por_via_4cut  por_via_4cut_3
timestamp 1718283729
transform -1 0 20299 0 -1 -300491
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_18
timestamp 1718283729
transform 0 -1 9676 1 0 -305162
box 15948 -7932 16222 -7868
use comparator_final  x1
timestamp 1721068816
transform 1 0 6296 0 1 -286728
box -1988 -5804 11208 -1484
use delayPulse_final  x2
timestamp 1721073345
transform 1 0 1048 0 1 -2959
box 1311 -297437 38614 -274935
use sky130_fd_pr__nfet_05v0_nvt_CZFQWY  XM2 paramcells
timestamp 1718283729
transform 1 0 15668 0 1 -288416
box -318 -567 318 567
use sky130_fd_pr__res_xhigh_po_0p35_NZA8SD  XR1 paramcells
timestamp 1718283729
transform -1 0 9633 0 1 -287413
box -2193 -1582 2193 1582
use sky130_fd_pr__res_xhigh_po_0p35_D2SRCG  XR10 paramcells
timestamp 1718283729
transform -1 0 12161 0 1 -287431
box -201 -1482 201 1482
use sky130_fd_pr__res_xhigh_po_0p35_SZAJAG  XR12 paramcells
timestamp 1718283729
transform -1 0 13843 0 1 -287413
box -1363 -1582 1363 1582
<< labels >>
flabel metal2 39385 -287337 39585 -287137 0 FreeSans 256 0 0 0 porb_h
port 7 nsew
flabel metal2 39296 -289388 39496 -289188 0 FreeSans 256 0 0 0 porb
port 5 nsew
flabel metal2 39301 -290929 39501 -290729 0 FreeSans 256 0 0 0 por
port 1 nsew
flabel metal2 24555 -293294 24755 -293094 0 FreeSans 256 0 0 0 dvss
port 6 nsew
flabel metal2 39292 -290256 39492 -290056 0 FreeSans 256 0 0 0 dvdd
port 4 nsew
flabel metal2 3491 -289455 3691 -289255 0 FreeSans 256 0 0 0 avdd
port 3 nsew
flabel metal2 3569 -292649 3769 -292449 0 FreeSans 256 0 0 0 vbg
port 0 nsew
flabel metal2 3612 -293264 3812 -293064 0 FreeSans 256 0 0 0 avss
port 2 nsew
<< end >>
