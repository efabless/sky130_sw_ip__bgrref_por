magic
tech sky130A
magscale 1 2
timestamp 1717613630
<< error_p >>
rect -29 472 29 478
rect -29 438 -17 472
rect -29 432 29 438
rect -29 -438 29 -432
rect -29 -472 -17 -438
rect -29 -478 29 -472
<< pwell >>
rect -226 -610 226 610
<< nmos >>
rect -30 -400 30 400
<< ndiff >>
rect -88 388 -30 400
rect -88 -388 -76 388
rect -42 -388 -30 388
rect -88 -400 -30 -388
rect 30 388 88 400
rect 30 -388 42 388
rect 76 -388 88 388
rect 30 -400 88 -388
<< ndiffc >>
rect -76 -388 -42 388
rect 42 -388 76 388
<< psubdiff >>
rect -190 540 -94 574
rect 94 540 190 574
rect -190 478 -156 540
rect 156 478 190 540
rect -190 -540 -156 -478
rect 156 -540 190 -478
rect -190 -574 -94 -540
rect 94 -574 190 -540
<< psubdiffcont >>
rect -94 540 94 574
rect -190 -478 -156 478
rect 156 -478 190 478
rect -94 -574 94 -540
<< poly >>
rect -33 472 33 488
rect -33 438 -17 472
rect 17 438 33 472
rect -33 422 33 438
rect -30 400 30 422
rect -30 -422 30 -400
rect -33 -438 33 -422
rect -33 -472 -17 -438
rect 17 -472 33 -438
rect -33 -488 33 -472
<< polycont >>
rect -17 438 17 472
rect -17 -472 17 -438
<< locali >>
rect -190 540 -94 574
rect 94 540 190 574
rect -190 478 -156 540
rect 156 478 190 540
rect -33 438 -17 472
rect 17 438 33 472
rect -76 388 -42 404
rect -76 -404 -42 -388
rect 42 388 76 404
rect 42 -404 76 -388
rect -33 -472 -17 -438
rect 17 -472 33 -438
rect -190 -540 -156 -478
rect 156 -540 190 -478
rect -190 -574 -94 -540
rect 94 -574 190 -540
<< viali >>
rect -17 438 17 472
rect -76 -388 -42 388
rect 42 -388 76 388
rect -17 -472 17 -438
<< metal1 >>
rect -29 472 29 478
rect -29 438 -17 472
rect 17 438 29 472
rect -29 432 29 438
rect -82 388 -36 400
rect -82 -388 -76 388
rect -42 -388 -36 388
rect -82 -400 -36 -388
rect 36 388 82 400
rect 36 -388 42 388
rect 76 -388 82 388
rect 36 -400 82 -388
rect -29 -438 29 -432
rect -29 -472 -17 -438
rect 17 -472 29 -438
rect -29 -478 29 -472
<< properties >>
string FIXED_BBOX -173 -557 173 557
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4.0 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
