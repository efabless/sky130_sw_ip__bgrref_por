magic
tech sky130A
magscale 1 2
timestamp 1717363523
<< pwell >>
rect -201 -25582 201 25582
<< psubdiff >>
rect -165 25512 -69 25546
rect 69 25512 165 25546
rect -165 25450 -131 25512
rect 131 25450 165 25512
rect -165 -25512 -131 -25450
rect 131 -25512 165 -25450
rect -165 -25546 -69 -25512
rect 69 -25546 165 -25512
<< psubdiffcont >>
rect -69 25512 69 25546
rect -165 -25450 -131 25450
rect 131 -25450 165 25450
rect -69 -25546 69 -25512
<< xpolycontact >>
rect -35 24984 35 25416
rect -35 -25416 35 -24984
<< xpolyres >>
rect -35 -24984 35 24984
<< locali >>
rect -165 25512 -69 25546
rect 69 25512 165 25546
rect -165 25450 -131 25512
rect 131 25450 165 25512
rect -165 -25512 -131 -25450
rect 131 -25512 165 -25450
rect -165 -25546 -69 -25512
rect 69 -25546 165 -25512
<< viali >>
rect -19 25001 19 25398
rect -19 -25398 19 -25001
<< metal1 >>
rect -25 25398 25 25410
rect -25 25001 -19 25398
rect 19 25001 25 25398
rect -25 24989 25 25001
rect -25 -25001 25 -24989
rect -25 -25398 -19 -25001
rect 19 -25398 25 -25001
rect -25 -25410 25 -25398
<< properties >>
string FIXED_BBOX -148 -25529 148 25529
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 250.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 1.429meg dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
