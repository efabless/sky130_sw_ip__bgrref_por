magic
tech sky130A
timestamp 1717527227
<< metal1 >>
rect 8044 -3963 8047 -3937
rect 8108 -3963 8111 -3937
<< via1 >>
rect 8047 -3963 8108 -3937
<< metal2 >>
rect 8047 -3937 8108 -3934
rect 8047 -3966 8108 -3963
<< end >>
