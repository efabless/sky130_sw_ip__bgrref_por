magic
tech sky130A
magscale 1 2
timestamp 1718283729
<< metal4 >>
rect -4098 17839 -200 17880
rect -4098 14561 -456 17839
rect -220 14561 -200 17839
rect -4098 14520 -200 14561
rect 200 17839 4098 17880
rect 200 14561 3842 17839
rect 4078 14561 4098 17839
rect 200 14520 4098 14561
rect -4098 14239 -200 14280
rect -4098 10961 -456 14239
rect -220 10961 -200 14239
rect -4098 10920 -200 10961
rect 200 14239 4098 14280
rect 200 10961 3842 14239
rect 4078 10961 4098 14239
rect 200 10920 4098 10961
rect -4098 10639 -200 10680
rect -4098 7361 -456 10639
rect -220 7361 -200 10639
rect -4098 7320 -200 7361
rect 200 10639 4098 10680
rect 200 7361 3842 10639
rect 4078 7361 4098 10639
rect 200 7320 4098 7361
rect -4098 7039 -200 7080
rect -4098 3761 -456 7039
rect -220 3761 -200 7039
rect -4098 3720 -200 3761
rect 200 7039 4098 7080
rect 200 3761 3842 7039
rect 4078 3761 4098 7039
rect 200 3720 4098 3761
rect -4098 3439 -200 3480
rect -4098 161 -456 3439
rect -220 161 -200 3439
rect -4098 120 -200 161
rect 200 3439 4098 3480
rect 200 161 3842 3439
rect 4078 161 4098 3439
rect 200 120 4098 161
rect -4098 -161 -200 -120
rect -4098 -3439 -456 -161
rect -220 -3439 -200 -161
rect -4098 -3480 -200 -3439
rect 200 -161 4098 -120
rect 200 -3439 3842 -161
rect 4078 -3439 4098 -161
rect 200 -3480 4098 -3439
rect -4098 -3761 -200 -3720
rect -4098 -7039 -456 -3761
rect -220 -7039 -200 -3761
rect -4098 -7080 -200 -7039
rect 200 -3761 4098 -3720
rect 200 -7039 3842 -3761
rect 4078 -7039 4098 -3761
rect 200 -7080 4098 -7039
rect -4098 -7361 -200 -7320
rect -4098 -10639 -456 -7361
rect -220 -10639 -200 -7361
rect -4098 -10680 -200 -10639
rect 200 -7361 4098 -7320
rect 200 -10639 3842 -7361
rect 4078 -10639 4098 -7361
rect 200 -10680 4098 -10639
rect -4098 -10961 -200 -10920
rect -4098 -14239 -456 -10961
rect -220 -14239 -200 -10961
rect -4098 -14280 -200 -14239
rect 200 -10961 4098 -10920
rect 200 -14239 3842 -10961
rect 4078 -14239 4098 -10961
rect 200 -14280 4098 -14239
rect -4098 -14561 -200 -14520
rect -4098 -17839 -456 -14561
rect -220 -17839 -200 -14561
rect -4098 -17880 -200 -17839
rect 200 -14561 4098 -14520
rect 200 -17839 3842 -14561
rect 4078 -17839 4098 -14561
rect 200 -17880 4098 -17839
<< via4 >>
rect -456 14561 -220 17839
rect 3842 14561 4078 17839
rect -456 10961 -220 14239
rect 3842 10961 4078 14239
rect -456 7361 -220 10639
rect 3842 7361 4078 10639
rect -456 3761 -220 7039
rect 3842 3761 4078 7039
rect -456 161 -220 3439
rect 3842 161 4078 3439
rect -456 -3439 -220 -161
rect 3842 -3439 4078 -161
rect -456 -7039 -220 -3761
rect 3842 -7039 4078 -3761
rect -456 -10639 -220 -7361
rect 3842 -10639 4078 -7361
rect -456 -14239 -220 -10961
rect 3842 -14239 4078 -10961
rect -456 -17839 -220 -14561
rect 3842 -17839 4078 -14561
<< mimcap2 >>
rect -4018 17760 -818 17800
rect -4018 14640 -3978 17760
rect -858 14640 -818 17760
rect -4018 14600 -818 14640
rect 280 17760 3480 17800
rect 280 14640 320 17760
rect 3440 14640 3480 17760
rect 280 14600 3480 14640
rect -4018 14160 -818 14200
rect -4018 11040 -3978 14160
rect -858 11040 -818 14160
rect -4018 11000 -818 11040
rect 280 14160 3480 14200
rect 280 11040 320 14160
rect 3440 11040 3480 14160
rect 280 11000 3480 11040
rect -4018 10560 -818 10600
rect -4018 7440 -3978 10560
rect -858 7440 -818 10560
rect -4018 7400 -818 7440
rect 280 10560 3480 10600
rect 280 7440 320 10560
rect 3440 7440 3480 10560
rect 280 7400 3480 7440
rect -4018 6960 -818 7000
rect -4018 3840 -3978 6960
rect -858 3840 -818 6960
rect -4018 3800 -818 3840
rect 280 6960 3480 7000
rect 280 3840 320 6960
rect 3440 3840 3480 6960
rect 280 3800 3480 3840
rect -4018 3360 -818 3400
rect -4018 240 -3978 3360
rect -858 240 -818 3360
rect -4018 200 -818 240
rect 280 3360 3480 3400
rect 280 240 320 3360
rect 3440 240 3480 3360
rect 280 200 3480 240
rect -4018 -240 -818 -200
rect -4018 -3360 -3978 -240
rect -858 -3360 -818 -240
rect -4018 -3400 -818 -3360
rect 280 -240 3480 -200
rect 280 -3360 320 -240
rect 3440 -3360 3480 -240
rect 280 -3400 3480 -3360
rect -4018 -3840 -818 -3800
rect -4018 -6960 -3978 -3840
rect -858 -6960 -818 -3840
rect -4018 -7000 -818 -6960
rect 280 -3840 3480 -3800
rect 280 -6960 320 -3840
rect 3440 -6960 3480 -3840
rect 280 -7000 3480 -6960
rect -4018 -7440 -818 -7400
rect -4018 -10560 -3978 -7440
rect -858 -10560 -818 -7440
rect -4018 -10600 -818 -10560
rect 280 -7440 3480 -7400
rect 280 -10560 320 -7440
rect 3440 -10560 3480 -7440
rect 280 -10600 3480 -10560
rect -4018 -11040 -818 -11000
rect -4018 -14160 -3978 -11040
rect -858 -14160 -818 -11040
rect -4018 -14200 -818 -14160
rect 280 -11040 3480 -11000
rect 280 -14160 320 -11040
rect 3440 -14160 3480 -11040
rect 280 -14200 3480 -14160
rect -4018 -14640 -818 -14600
rect -4018 -17760 -3978 -14640
rect -858 -17760 -818 -14640
rect -4018 -17800 -818 -17760
rect 280 -14640 3480 -14600
rect 280 -17760 320 -14640
rect 3440 -17760 3480 -14640
rect 280 -17800 3480 -17760
<< mimcap2contact >>
rect -3978 14640 -858 17760
rect 320 14640 3440 17760
rect -3978 11040 -858 14160
rect 320 11040 3440 14160
rect -3978 7440 -858 10560
rect 320 7440 3440 10560
rect -3978 3840 -858 6960
rect 320 3840 3440 6960
rect -3978 240 -858 3360
rect 320 240 3440 3360
rect -3978 -3360 -858 -240
rect 320 -3360 3440 -240
rect -3978 -6960 -858 -3840
rect 320 -6960 3440 -3840
rect -3978 -10560 -858 -7440
rect 320 -10560 3440 -7440
rect -3978 -14160 -858 -11040
rect 320 -14160 3440 -11040
rect -3978 -17760 -858 -14640
rect 320 -17760 3440 -14640
<< metal5 >>
rect -2578 17784 -2258 18000
rect -498 17839 -178 18000
rect -4002 17760 -834 17784
rect -4002 14640 -3978 17760
rect -858 14640 -834 17760
rect -4002 14616 -834 14640
rect -2578 14184 -2258 14616
rect -498 14561 -456 17839
rect -220 14561 -178 17839
rect 1720 17784 2040 18000
rect 3800 17839 4120 18000
rect 296 17760 3464 17784
rect 296 14640 320 17760
rect 3440 14640 3464 17760
rect 296 14616 3464 14640
rect -498 14239 -178 14561
rect -4002 14160 -834 14184
rect -4002 11040 -3978 14160
rect -858 11040 -834 14160
rect -4002 11016 -834 11040
rect -2578 10584 -2258 11016
rect -498 10961 -456 14239
rect -220 10961 -178 14239
rect 1720 14184 2040 14616
rect 3800 14561 3842 17839
rect 4078 14561 4120 17839
rect 3800 14239 4120 14561
rect 296 14160 3464 14184
rect 296 11040 320 14160
rect 3440 11040 3464 14160
rect 296 11016 3464 11040
rect -498 10639 -178 10961
rect -4002 10560 -834 10584
rect -4002 7440 -3978 10560
rect -858 7440 -834 10560
rect -4002 7416 -834 7440
rect -2578 6984 -2258 7416
rect -498 7361 -456 10639
rect -220 7361 -178 10639
rect 1720 10584 2040 11016
rect 3800 10961 3842 14239
rect 4078 10961 4120 14239
rect 3800 10639 4120 10961
rect 296 10560 3464 10584
rect 296 7440 320 10560
rect 3440 7440 3464 10560
rect 296 7416 3464 7440
rect -498 7039 -178 7361
rect -4002 6960 -834 6984
rect -4002 3840 -3978 6960
rect -858 3840 -834 6960
rect -4002 3816 -834 3840
rect -2578 3384 -2258 3816
rect -498 3761 -456 7039
rect -220 3761 -178 7039
rect 1720 6984 2040 7416
rect 3800 7361 3842 10639
rect 4078 7361 4120 10639
rect 3800 7039 4120 7361
rect 296 6960 3464 6984
rect 296 3840 320 6960
rect 3440 3840 3464 6960
rect 296 3816 3464 3840
rect -498 3439 -178 3761
rect -4002 3360 -834 3384
rect -4002 240 -3978 3360
rect -858 240 -834 3360
rect -4002 216 -834 240
rect -2578 -216 -2258 216
rect -498 161 -456 3439
rect -220 161 -178 3439
rect 1720 3384 2040 3816
rect 3800 3761 3842 7039
rect 4078 3761 4120 7039
rect 3800 3439 4120 3761
rect 296 3360 3464 3384
rect 296 240 320 3360
rect 3440 240 3464 3360
rect 296 216 3464 240
rect -498 -161 -178 161
rect -4002 -240 -834 -216
rect -4002 -3360 -3978 -240
rect -858 -3360 -834 -240
rect -4002 -3384 -834 -3360
rect -2578 -3816 -2258 -3384
rect -498 -3439 -456 -161
rect -220 -3439 -178 -161
rect 1720 -216 2040 216
rect 3800 161 3842 3439
rect 4078 161 4120 3439
rect 3800 -161 4120 161
rect 296 -240 3464 -216
rect 296 -3360 320 -240
rect 3440 -3360 3464 -240
rect 296 -3384 3464 -3360
rect -498 -3761 -178 -3439
rect -4002 -3840 -834 -3816
rect -4002 -6960 -3978 -3840
rect -858 -6960 -834 -3840
rect -4002 -6984 -834 -6960
rect -2578 -7416 -2258 -6984
rect -498 -7039 -456 -3761
rect -220 -7039 -178 -3761
rect 1720 -3816 2040 -3384
rect 3800 -3439 3842 -161
rect 4078 -3439 4120 -161
rect 3800 -3761 4120 -3439
rect 296 -3840 3464 -3816
rect 296 -6960 320 -3840
rect 3440 -6960 3464 -3840
rect 296 -6984 3464 -6960
rect -498 -7361 -178 -7039
rect -4002 -7440 -834 -7416
rect -4002 -10560 -3978 -7440
rect -858 -10560 -834 -7440
rect -4002 -10584 -834 -10560
rect -2578 -11016 -2258 -10584
rect -498 -10639 -456 -7361
rect -220 -10639 -178 -7361
rect 1720 -7416 2040 -6984
rect 3800 -7039 3842 -3761
rect 4078 -7039 4120 -3761
rect 3800 -7361 4120 -7039
rect 296 -7440 3464 -7416
rect 296 -10560 320 -7440
rect 3440 -10560 3464 -7440
rect 296 -10584 3464 -10560
rect -498 -10961 -178 -10639
rect -4002 -11040 -834 -11016
rect -4002 -14160 -3978 -11040
rect -858 -14160 -834 -11040
rect -4002 -14184 -834 -14160
rect -2578 -14616 -2258 -14184
rect -498 -14239 -456 -10961
rect -220 -14239 -178 -10961
rect 1720 -11016 2040 -10584
rect 3800 -10639 3842 -7361
rect 4078 -10639 4120 -7361
rect 3800 -10961 4120 -10639
rect 296 -11040 3464 -11016
rect 296 -14160 320 -11040
rect 3440 -14160 3464 -11040
rect 296 -14184 3464 -14160
rect -498 -14561 -178 -14239
rect -4002 -14640 -834 -14616
rect -4002 -17760 -3978 -14640
rect -858 -17760 -834 -14640
rect -4002 -17784 -834 -17760
rect -2578 -18000 -2258 -17784
rect -498 -17839 -456 -14561
rect -220 -17839 -178 -14561
rect 1720 -14616 2040 -14184
rect 3800 -14239 3842 -10961
rect 4078 -14239 4120 -10961
rect 3800 -14561 4120 -14239
rect 296 -14640 3464 -14616
rect 296 -17760 320 -14640
rect 3440 -17760 3464 -14640
rect 296 -17784 3464 -17760
rect -498 -18000 -178 -17839
rect 1720 -18000 2040 -17784
rect 3800 -17839 3842 -14561
rect 4078 -17839 4120 -14561
rect 3800 -18000 4120 -17839
<< properties >>
string FIXED_BBOX 200 14520 3560 17880
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 16.0 l 16.0 val 524.159 carea 2.00 cperi 0.19 nx 2 ny 10 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
