magic
tech sky130A
magscale 1 2
timestamp 1717528722
<< metal3 >>
rect -4192 18954 -720 18982
rect -4192 15930 -804 18954
rect -740 15930 -720 18954
rect -4192 15902 -720 15930
rect 120 18954 3592 18982
rect 120 15930 3508 18954
rect 3572 15930 3592 18954
rect 120 15902 3592 15930
rect -4192 15356 -720 15384
rect -4192 12332 -804 15356
rect -740 12332 -720 15356
rect -4192 12304 -720 12332
rect 120 15356 3592 15384
rect 120 12332 3508 15356
rect 3572 12332 3592 15356
rect 120 12304 3592 12332
rect -4192 11758 -720 11786
rect -4192 8734 -804 11758
rect -740 8734 -720 11758
rect -4192 8706 -720 8734
rect 120 11758 3592 11786
rect 120 8734 3508 11758
rect 3572 8734 3592 11758
rect 120 8706 3592 8734
rect -4192 8160 -720 8188
rect -4192 5136 -804 8160
rect -740 5136 -720 8160
rect -4192 5108 -720 5136
rect 120 8160 3592 8188
rect 120 5136 3508 8160
rect 3572 5136 3592 8160
rect 120 5108 3592 5136
rect -4192 4562 -720 4590
rect -4192 1538 -804 4562
rect -740 1538 -720 4562
rect -4192 1510 -720 1538
rect 120 4562 3592 4590
rect 120 1538 3508 4562
rect 3572 1538 3592 4562
rect 120 1510 3592 1538
rect -4192 964 -720 992
rect -4192 -2060 -804 964
rect -740 -2060 -720 964
rect -4192 -2088 -720 -2060
rect 120 964 3592 992
rect 120 -2060 3508 964
rect 3572 -2060 3592 964
rect 120 -2088 3592 -2060
rect -4192 -2634 -720 -2606
rect -4192 -5658 -804 -2634
rect -740 -5658 -720 -2634
rect -4192 -5686 -720 -5658
rect 120 -2634 3592 -2606
rect 120 -5658 3508 -2634
rect 3572 -5658 3592 -2634
rect 120 -5686 3592 -5658
rect -4192 -6232 -720 -6204
rect -4192 -9256 -804 -6232
rect -740 -9256 -720 -6232
rect -4192 -9284 -720 -9256
rect 120 -6232 3592 -6204
rect 120 -9256 3508 -6232
rect 3572 -9256 3592 -6232
rect 120 -9284 3592 -9256
rect -4192 -9830 -720 -9802
rect -4192 -12854 -804 -9830
rect -740 -12854 -720 -9830
rect -4192 -12882 -720 -12854
rect 120 -9830 3592 -9802
rect 120 -12854 3508 -9830
rect 3572 -12854 3592 -9830
rect 120 -12882 3592 -12854
rect -4192 -13428 -720 -13400
rect -4192 -16452 -804 -13428
rect -740 -16452 -720 -13428
rect -4192 -16480 -720 -16452
rect 120 -13428 3592 -13400
rect 120 -16452 3508 -13428
rect 3572 -16452 3592 -13428
rect 120 -16480 3592 -16452
<< via3 >>
rect -804 15930 -740 18954
rect 3508 15930 3572 18954
rect -804 12332 -740 15356
rect 3508 12332 3572 15356
rect -804 8734 -740 11758
rect 3508 8734 3572 11758
rect -804 5136 -740 8160
rect 3508 5136 3572 8160
rect -804 1538 -740 4562
rect 3508 1538 3572 4562
rect -804 -2060 -740 964
rect 3508 -2060 3572 964
rect -804 -5658 -740 -2634
rect 3508 -5658 3572 -2634
rect -804 -9256 -740 -6232
rect 3508 -9256 3572 -6232
rect -804 -12854 -740 -9830
rect 3508 -12854 3572 -9830
rect -804 -16452 -740 -13428
rect 3508 -16452 3572 -13428
<< mimcap >>
rect -4152 18902 -1152 18942
rect -4152 15982 -4112 18902
rect -1192 15982 -1152 18902
rect -4152 15942 -1152 15982
rect 160 18902 3160 18942
rect 160 15982 200 18902
rect 3120 15982 3160 18902
rect 160 15942 3160 15982
rect -4152 15304 -1152 15344
rect -4152 12384 -4112 15304
rect -1192 12384 -1152 15304
rect -4152 12344 -1152 12384
rect 160 15304 3160 15344
rect 160 12384 200 15304
rect 3120 12384 3160 15304
rect 160 12344 3160 12384
rect -4152 11706 -1152 11746
rect -4152 8786 -4112 11706
rect -1192 8786 -1152 11706
rect -4152 8746 -1152 8786
rect 160 11706 3160 11746
rect 160 8786 200 11706
rect 3120 8786 3160 11706
rect 160 8746 3160 8786
rect -4152 8108 -1152 8148
rect -4152 5188 -4112 8108
rect -1192 5188 -1152 8108
rect -4152 5148 -1152 5188
rect 160 8108 3160 8148
rect 160 5188 200 8108
rect 3120 5188 3160 8108
rect 160 5148 3160 5188
rect -4152 4510 -1152 4550
rect -4152 1590 -4112 4510
rect -1192 1590 -1152 4510
rect -4152 1550 -1152 1590
rect 160 4510 3160 4550
rect 160 1590 200 4510
rect 3120 1590 3160 4510
rect 160 1550 3160 1590
rect -4152 912 -1152 952
rect -4152 -2008 -4112 912
rect -1192 -2008 -1152 912
rect -4152 -2048 -1152 -2008
rect 160 912 3160 952
rect 160 -2008 200 912
rect 3120 -2008 3160 912
rect 160 -2048 3160 -2008
rect -4152 -2686 -1152 -2646
rect -4152 -5606 -4112 -2686
rect -1192 -5606 -1152 -2686
rect -4152 -5646 -1152 -5606
rect 160 -2686 3160 -2646
rect 160 -5606 200 -2686
rect 3120 -5606 3160 -2686
rect 160 -5646 3160 -5606
rect -4152 -6284 -1152 -6244
rect -4152 -9204 -4112 -6284
rect -1192 -9204 -1152 -6284
rect -4152 -9244 -1152 -9204
rect 160 -6284 3160 -6244
rect 160 -9204 200 -6284
rect 3120 -9204 3160 -6284
rect 160 -9244 3160 -9204
rect -4152 -9882 -1152 -9842
rect -4152 -12802 -4112 -9882
rect -1192 -12802 -1152 -9882
rect -4152 -12842 -1152 -12802
rect 160 -9882 3160 -9842
rect 160 -12802 200 -9882
rect 3120 -12802 3160 -9882
rect 160 -12842 3160 -12802
rect -4152 -13480 -1152 -13440
rect -4152 -16400 -4112 -13480
rect -1192 -16400 -1152 -13480
rect -4152 -16440 -1152 -16400
rect 160 -13480 3160 -13440
rect 160 -16400 200 -13480
rect 3120 -16400 3160 -13480
rect 160 -16440 3160 -16400
<< mimcapcontact >>
rect -4112 15982 -1192 18902
rect 200 15982 3120 18902
rect -4112 12384 -1192 15304
rect 200 12384 3120 15304
rect -4112 8786 -1192 11706
rect 200 8786 3120 11706
rect -4112 5188 -1192 8108
rect 200 5188 3120 8108
rect -4112 1590 -1192 4510
rect 200 1590 3120 4510
rect -4112 -2008 -1192 912
rect 200 -2008 3120 912
rect -4112 -5606 -1192 -2686
rect 200 -5606 3120 -2686
rect -4112 -9204 -1192 -6284
rect 200 -9204 3120 -6284
rect -4112 -12802 -1192 -9882
rect 200 -12802 3120 -9882
rect -4112 -16400 -1192 -13480
rect 200 -16400 3120 -13480
<< metal4 >>
rect -2704 18903 -2600 19102
rect -824 18954 -720 19102
rect -4113 18902 -1191 18903
rect -4113 15982 -4112 18902
rect -1192 15982 -1191 18902
rect -4113 15981 -1191 15982
rect -2704 15305 -2600 15981
rect -824 15930 -804 18954
rect -740 15930 -720 18954
rect 1608 18903 1712 19102
rect 3488 18954 3592 19102
rect 199 18902 3121 18903
rect 199 15982 200 18902
rect 3120 15982 3121 18902
rect 199 15981 3121 15982
rect -824 15356 -720 15930
rect -4113 15304 -1191 15305
rect -4113 12384 -4112 15304
rect -1192 12384 -1191 15304
rect -4113 12383 -1191 12384
rect -2704 11707 -2600 12383
rect -824 12332 -804 15356
rect -740 12332 -720 15356
rect 1608 15305 1712 15981
rect 3488 15930 3508 18954
rect 3572 15930 3592 18954
rect 3488 15356 3592 15930
rect 199 15304 3121 15305
rect 199 12384 200 15304
rect 3120 12384 3121 15304
rect 199 12383 3121 12384
rect -824 11758 -720 12332
rect -4113 11706 -1191 11707
rect -4113 8786 -4112 11706
rect -1192 8786 -1191 11706
rect -4113 8785 -1191 8786
rect -2704 8109 -2600 8785
rect -824 8734 -804 11758
rect -740 8734 -720 11758
rect 1608 11707 1712 12383
rect 3488 12332 3508 15356
rect 3572 12332 3592 15356
rect 3488 11758 3592 12332
rect 199 11706 3121 11707
rect 199 8786 200 11706
rect 3120 8786 3121 11706
rect 199 8785 3121 8786
rect -824 8160 -720 8734
rect -4113 8108 -1191 8109
rect -4113 5188 -4112 8108
rect -1192 5188 -1191 8108
rect -4113 5187 -1191 5188
rect -2704 4511 -2600 5187
rect -824 5136 -804 8160
rect -740 5136 -720 8160
rect 1608 8109 1712 8785
rect 3488 8734 3508 11758
rect 3572 8734 3592 11758
rect 3488 8160 3592 8734
rect 199 8108 3121 8109
rect 199 5188 200 8108
rect 3120 5188 3121 8108
rect 199 5187 3121 5188
rect -824 4562 -720 5136
rect -4113 4510 -1191 4511
rect -4113 1590 -4112 4510
rect -1192 1590 -1191 4510
rect -4113 1589 -1191 1590
rect -2704 913 -2600 1589
rect -824 1538 -804 4562
rect -740 1538 -720 4562
rect 1608 4511 1712 5187
rect 3488 5136 3508 8160
rect 3572 5136 3592 8160
rect 3488 4562 3592 5136
rect 199 4510 3121 4511
rect 199 1590 200 4510
rect 3120 1590 3121 4510
rect 199 1589 3121 1590
rect -824 964 -720 1538
rect -4113 912 -1191 913
rect -4113 -2008 -4112 912
rect -1192 -2008 -1191 912
rect -4113 -2009 -1191 -2008
rect -2704 -2685 -2600 -2009
rect -824 -2060 -804 964
rect -740 -2060 -720 964
rect 1608 913 1712 1589
rect 3488 1538 3508 4562
rect 3572 1538 3592 4562
rect 3488 964 3592 1538
rect 199 912 3121 913
rect 199 -2008 200 912
rect 3120 -2008 3121 912
rect 199 -2009 3121 -2008
rect -824 -2634 -720 -2060
rect -4113 -2686 -1191 -2685
rect -4113 -5606 -4112 -2686
rect -1192 -5606 -1191 -2686
rect -4113 -5607 -1191 -5606
rect -2704 -6283 -2600 -5607
rect -824 -5658 -804 -2634
rect -740 -5658 -720 -2634
rect 1608 -2685 1712 -2009
rect 3488 -2060 3508 964
rect 3572 -2060 3592 964
rect 3488 -2634 3592 -2060
rect 199 -2686 3121 -2685
rect 199 -5606 200 -2686
rect 3120 -5606 3121 -2686
rect 199 -5607 3121 -5606
rect -824 -6232 -720 -5658
rect -4113 -6284 -1191 -6283
rect -4113 -9204 -4112 -6284
rect -1192 -9204 -1191 -6284
rect -4113 -9205 -1191 -9204
rect -2704 -9881 -2600 -9205
rect -824 -9256 -804 -6232
rect -740 -9256 -720 -6232
rect 1608 -6283 1712 -5607
rect 3488 -5658 3508 -2634
rect 3572 -5658 3592 -2634
rect 3488 -6232 3592 -5658
rect 199 -6284 3121 -6283
rect 199 -9204 200 -6284
rect 3120 -9204 3121 -6284
rect 199 -9205 3121 -9204
rect -824 -9830 -720 -9256
rect -4113 -9882 -1191 -9881
rect -4113 -12802 -4112 -9882
rect -1192 -12802 -1191 -9882
rect -4113 -12803 -1191 -12802
rect -2704 -13479 -2600 -12803
rect -824 -12854 -804 -9830
rect -740 -12854 -720 -9830
rect 1608 -9881 1712 -9205
rect 3488 -9256 3508 -6232
rect 3572 -9256 3592 -6232
rect 3488 -9830 3592 -9256
rect 199 -9882 3121 -9881
rect 199 -12802 200 -9882
rect 3120 -12802 3121 -9882
rect 199 -12803 3121 -12802
rect -824 -13428 -720 -12854
rect -4113 -13480 -1191 -13479
rect -4113 -16400 -4112 -13480
rect -1192 -16400 -1191 -13480
rect -4113 -16401 -1191 -16400
rect -2704 -16600 -2600 -16401
rect -824 -16452 -804 -13428
rect -740 -16452 -720 -13428
rect 1608 -13479 1712 -12803
rect 3488 -12854 3508 -9830
rect 3572 -12854 3592 -9830
rect 3488 -13428 3592 -12854
rect 199 -13480 3121 -13479
rect 199 -16400 200 -13480
rect 3120 -16400 3121 -13480
rect 199 -16401 3121 -16400
rect -824 -16600 -720 -16452
rect 1608 -16600 1712 -16401
rect 3488 -16452 3508 -13428
rect 3572 -16452 3592 -13428
rect 3488 -16600 3592 -16452
<< properties >>
string FIXED_BBOX 120 13400 3200 16480
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 15.00 l 15.00 val 461.4 carea 2.00 cperi 0.19 nx 2 ny 10 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
