magic
tech sky130A
magscale 1 2
timestamp 1717527227
<< nwell >>
rect -387 -547 387 547
<< mvpmos >>
rect -129 -250 -29 250
rect 29 -250 129 250
<< mvpdiff >>
rect -187 238 -129 250
rect -187 -238 -175 238
rect -141 -238 -129 238
rect -187 -250 -129 -238
rect -29 238 29 250
rect -29 -238 -17 238
rect 17 -238 29 238
rect -29 -250 29 -238
rect 129 238 187 250
rect 129 -238 141 238
rect 175 -238 187 238
rect 129 -250 187 -238
<< mvpdiffc >>
rect -175 -238 -141 238
rect -17 -238 17 238
rect 141 -238 175 238
<< mvnsubdiff >>
rect -321 469 321 481
rect -321 435 -213 469
rect 213 435 321 469
rect -321 423 321 435
rect -321 373 -263 423
rect -321 -373 -309 373
rect -275 -373 -263 373
rect 263 373 321 423
rect -321 -423 -263 -373
rect 263 -373 275 373
rect 309 -373 321 373
rect 263 -423 321 -373
rect -321 -435 321 -423
rect -321 -469 -213 -435
rect 213 -469 321 -435
rect -321 -481 321 -469
<< mvnsubdiffcont >>
rect -213 435 213 469
rect -309 -373 -275 373
rect 275 -373 309 373
rect -213 -469 213 -435
<< poly >>
rect -129 331 -29 347
rect -129 297 -113 331
rect -45 297 -29 331
rect -129 250 -29 297
rect 29 331 129 347
rect 29 297 45 331
rect 113 297 129 331
rect 29 250 129 297
rect -129 -297 -29 -250
rect -129 -331 -113 -297
rect -45 -331 -29 -297
rect -129 -347 -29 -331
rect 29 -297 129 -250
rect 29 -331 45 -297
rect 113 -331 129 -297
rect 29 -347 129 -331
<< polycont >>
rect -113 297 -45 331
rect 45 297 113 331
rect -113 -331 -45 -297
rect 45 -331 113 -297
<< locali >>
rect -309 435 -213 469
rect 213 435 309 469
rect -309 373 -275 435
rect 275 373 309 435
rect -129 297 -113 331
rect -45 297 -29 331
rect 29 297 45 331
rect 113 297 129 331
rect -175 238 -141 254
rect -175 -254 -141 -238
rect -17 238 17 254
rect -17 -254 17 -238
rect 141 238 175 254
rect 141 -254 175 -238
rect -129 -331 -113 -297
rect -45 -331 -29 -297
rect 29 -331 45 -297
rect 113 -331 129 -297
rect -309 -435 -275 -373
rect 275 -435 309 -373
rect -309 -469 -213 -435
rect 213 -469 309 -435
<< viali >>
rect -113 297 -45 331
rect 45 297 113 331
rect -175 -238 -141 238
rect -17 -238 17 238
rect 141 -238 175 238
rect -113 -331 -45 -297
rect 45 -331 113 -297
<< metal1 >>
rect -125 331 -33 337
rect -125 297 -113 331
rect -45 297 -33 331
rect -125 291 -33 297
rect 33 331 125 337
rect 33 297 45 331
rect 113 297 125 331
rect 33 291 125 297
rect -181 238 -135 250
rect -181 -238 -175 238
rect -141 -238 -135 238
rect -181 -250 -135 -238
rect -23 238 23 250
rect -23 -238 -17 238
rect 17 -238 23 238
rect -23 -250 23 -238
rect 135 238 181 250
rect 135 -238 141 238
rect 175 -238 181 238
rect 135 -250 181 -238
rect -125 -297 -33 -291
rect -125 -331 -113 -297
rect -45 -331 -33 -297
rect -125 -337 -33 -331
rect 33 -297 125 -291
rect 33 -331 45 -297
rect 113 -331 125 -297
rect 33 -337 125 -331
<< properties >>
string FIXED_BBOX -292 -452 292 452
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2.5 l 0.50 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
