magic
tech sky130A
magscale 1 2
timestamp 1717554641
<< metal3 >>
rect -4192 18154 -620 18182
rect -4192 14930 -704 18154
rect -640 14930 -620 18154
rect -4192 14902 -620 14930
rect 120 18154 3692 18182
rect 120 14930 3608 18154
rect 3672 14930 3692 18154
rect 120 14902 3692 14930
rect -4192 14556 -620 14584
rect -4192 11332 -704 14556
rect -640 11332 -620 14556
rect -4192 11304 -620 11332
rect 120 14556 3692 14584
rect 120 11332 3608 14556
rect 3672 11332 3692 14556
rect 120 11304 3692 11332
rect -4192 10958 -620 10986
rect -4192 7734 -704 10958
rect -640 7734 -620 10958
rect -4192 7706 -620 7734
rect 120 10958 3692 10986
rect 120 7734 3608 10958
rect 3672 7734 3692 10958
rect 120 7706 3692 7734
rect -4192 7360 -620 7388
rect -4192 4136 -704 7360
rect -640 4136 -620 7360
rect -4192 4108 -620 4136
rect 120 7360 3692 7388
rect 120 4136 3608 7360
rect 3672 4136 3692 7360
rect 120 4108 3692 4136
rect -4192 3762 -620 3790
rect -4192 538 -704 3762
rect -640 538 -620 3762
rect -4192 510 -620 538
rect 120 3762 3692 3790
rect 120 538 3608 3762
rect 3672 538 3692 3762
rect 120 510 3692 538
rect -4192 164 -620 192
rect -4192 -3060 -704 164
rect -640 -3060 -620 164
rect -4192 -3088 -620 -3060
rect 120 164 3692 192
rect 120 -3060 3608 164
rect 3672 -3060 3692 164
rect 120 -3088 3692 -3060
rect -4192 -3434 -620 -3406
rect -4192 -6658 -704 -3434
rect -640 -6658 -620 -3434
rect -4192 -6686 -620 -6658
rect 120 -3434 3692 -3406
rect 120 -6658 3608 -3434
rect 3672 -6658 3692 -3434
rect 120 -6686 3692 -6658
rect -4192 -7032 -620 -7004
rect -4192 -10256 -704 -7032
rect -640 -10256 -620 -7032
rect -4192 -10284 -620 -10256
rect 120 -7032 3692 -7004
rect 120 -10256 3608 -7032
rect 3672 -10256 3692 -7032
rect 120 -10284 3692 -10256
rect -4192 -10630 -620 -10602
rect -4192 -13854 -704 -10630
rect -640 -13854 -620 -10630
rect -4192 -13882 -620 -13854
rect 120 -10630 3692 -10602
rect 120 -13854 3608 -10630
rect 3672 -13854 3692 -10630
rect 120 -13882 3692 -13854
rect -4192 -14228 -620 -14200
rect -4192 -17452 -704 -14228
rect -640 -17452 -620 -14228
rect -4192 -17480 -620 -17452
rect 120 -14228 3692 -14200
rect 120 -17452 3608 -14228
rect 3672 -17452 3692 -14228
rect 120 -17480 3692 -17452
<< via3 >>
rect -704 14930 -640 18154
rect 3608 14930 3672 18154
rect -704 11332 -640 14556
rect 3608 11332 3672 14556
rect -704 7734 -640 10958
rect 3608 7734 3672 10958
rect -704 4136 -640 7360
rect 3608 4136 3672 7360
rect -704 538 -640 3762
rect 3608 538 3672 3762
rect -704 -3060 -640 164
rect 3608 -3060 3672 164
rect -704 -6658 -640 -3434
rect 3608 -6658 3672 -3434
rect -704 -10256 -640 -7032
rect 3608 -10256 3672 -7032
rect -704 -13854 -640 -10630
rect 3608 -13854 3672 -10630
rect -704 -17452 -640 -14228
rect 3608 -17452 3672 -14228
<< mimcap >>
rect -4152 18102 -952 18142
rect -4152 14982 -4112 18102
rect -992 14982 -952 18102
rect -4152 14942 -952 14982
rect 160 18102 3360 18142
rect 160 14982 200 18102
rect 3320 14982 3360 18102
rect 160 14942 3360 14982
rect -4152 14504 -952 14544
rect -4152 11384 -4112 14504
rect -992 11384 -952 14504
rect -4152 11344 -952 11384
rect 160 14504 3360 14544
rect 160 11384 200 14504
rect 3320 11384 3360 14504
rect 160 11344 3360 11384
rect -4152 10906 -952 10946
rect -4152 7786 -4112 10906
rect -992 7786 -952 10906
rect -4152 7746 -952 7786
rect 160 10906 3360 10946
rect 160 7786 200 10906
rect 3320 7786 3360 10906
rect 160 7746 3360 7786
rect -4152 7308 -952 7348
rect -4152 4188 -4112 7308
rect -992 4188 -952 7308
rect -4152 4148 -952 4188
rect 160 7308 3360 7348
rect 160 4188 200 7308
rect 3320 4188 3360 7308
rect 160 4148 3360 4188
rect -4152 3710 -952 3750
rect -4152 590 -4112 3710
rect -992 590 -952 3710
rect -4152 550 -952 590
rect 160 3710 3360 3750
rect 160 590 200 3710
rect 3320 590 3360 3710
rect 160 550 3360 590
rect -4152 112 -952 152
rect -4152 -3008 -4112 112
rect -992 -3008 -952 112
rect -4152 -3048 -952 -3008
rect 160 112 3360 152
rect 160 -3008 200 112
rect 3320 -3008 3360 112
rect 160 -3048 3360 -3008
rect -4152 -3486 -952 -3446
rect -4152 -6606 -4112 -3486
rect -992 -6606 -952 -3486
rect -4152 -6646 -952 -6606
rect 160 -3486 3360 -3446
rect 160 -6606 200 -3486
rect 3320 -6606 3360 -3486
rect 160 -6646 3360 -6606
rect -4152 -7084 -952 -7044
rect -4152 -10204 -4112 -7084
rect -992 -10204 -952 -7084
rect -4152 -10244 -952 -10204
rect 160 -7084 3360 -7044
rect 160 -10204 200 -7084
rect 3320 -10204 3360 -7084
rect 160 -10244 3360 -10204
rect -4152 -10682 -952 -10642
rect -4152 -13802 -4112 -10682
rect -992 -13802 -952 -10682
rect -4152 -13842 -952 -13802
rect 160 -10682 3360 -10642
rect 160 -13802 200 -10682
rect 3320 -13802 3360 -10682
rect 160 -13842 3360 -13802
rect -4152 -14280 -952 -14240
rect -4152 -17400 -4112 -14280
rect -992 -17400 -952 -14280
rect -4152 -17440 -952 -17400
rect 160 -14280 3360 -14240
rect 160 -17400 200 -14280
rect 3320 -17400 3360 -14280
rect 160 -17440 3360 -17400
<< mimcapcontact >>
rect -4112 14982 -992 18102
rect 200 14982 3320 18102
rect -4112 11384 -992 14504
rect 200 11384 3320 14504
rect -4112 7786 -992 10906
rect 200 7786 3320 10906
rect -4112 4188 -992 7308
rect 200 4188 3320 7308
rect -4112 590 -992 3710
rect 200 590 3320 3710
rect -4112 -3008 -992 112
rect 200 -3008 3320 112
rect -4112 -6606 -992 -3486
rect 200 -6606 3320 -3486
rect -4112 -10204 -992 -7084
rect 200 -10204 3320 -7084
rect -4112 -13802 -992 -10682
rect 200 -13802 3320 -10682
rect -4112 -17400 -992 -14280
rect 200 -17400 3320 -14280
<< metal4 >>
rect -2604 18103 -2500 18302
rect -724 18154 -620 18302
rect -4113 18102 -991 18103
rect -4113 14982 -4112 18102
rect -992 14982 -991 18102
rect -4113 14981 -991 14982
rect -2604 14505 -2500 14981
rect -724 14930 -704 18154
rect -640 14930 -620 18154
rect 1708 18103 1812 18302
rect 3588 18154 3692 18302
rect 199 18102 3321 18103
rect 199 14982 200 18102
rect 3320 14982 3321 18102
rect 199 14981 3321 14982
rect -724 14556 -620 14930
rect -4113 14504 -991 14505
rect -4113 11384 -4112 14504
rect -992 11384 -991 14504
rect -4113 11383 -991 11384
rect -2604 10907 -2500 11383
rect -724 11332 -704 14556
rect -640 11332 -620 14556
rect 1708 14505 1812 14981
rect 3588 14930 3608 18154
rect 3672 14930 3692 18154
rect 3588 14556 3692 14930
rect 199 14504 3321 14505
rect 199 11384 200 14504
rect 3320 11384 3321 14504
rect 199 11383 3321 11384
rect -724 10958 -620 11332
rect -4113 10906 -991 10907
rect -4113 7786 -4112 10906
rect -992 7786 -991 10906
rect -4113 7785 -991 7786
rect -2604 7309 -2500 7785
rect -724 7734 -704 10958
rect -640 7734 -620 10958
rect 1708 10907 1812 11383
rect 3588 11332 3608 14556
rect 3672 11332 3692 14556
rect 3588 10958 3692 11332
rect 199 10906 3321 10907
rect 199 7786 200 10906
rect 3320 7786 3321 10906
rect 199 7785 3321 7786
rect -724 7360 -620 7734
rect -4113 7308 -991 7309
rect -4113 4188 -4112 7308
rect -992 4188 -991 7308
rect -4113 4187 -991 4188
rect -2604 3711 -2500 4187
rect -724 4136 -704 7360
rect -640 4136 -620 7360
rect 1708 7309 1812 7785
rect 3588 7734 3608 10958
rect 3672 7734 3692 10958
rect 3588 7360 3692 7734
rect 199 7308 3321 7309
rect 199 4188 200 7308
rect 3320 4188 3321 7308
rect 199 4187 3321 4188
rect -724 3762 -620 4136
rect -4113 3710 -991 3711
rect -4113 590 -4112 3710
rect -992 590 -991 3710
rect -4113 589 -991 590
rect -2604 113 -2500 589
rect -724 538 -704 3762
rect -640 538 -620 3762
rect 1708 3711 1812 4187
rect 3588 4136 3608 7360
rect 3672 4136 3692 7360
rect 3588 3762 3692 4136
rect 199 3710 3321 3711
rect 199 590 200 3710
rect 3320 590 3321 3710
rect 199 589 3321 590
rect -724 164 -620 538
rect -4113 112 -991 113
rect -4113 -3008 -4112 112
rect -992 -3008 -991 112
rect -4113 -3009 -991 -3008
rect -2604 -3485 -2500 -3009
rect -724 -3060 -704 164
rect -640 -3060 -620 164
rect 1708 113 1812 589
rect 3588 538 3608 3762
rect 3672 538 3692 3762
rect 3588 164 3692 538
rect 199 112 3321 113
rect 199 -3008 200 112
rect 3320 -3008 3321 112
rect 199 -3009 3321 -3008
rect -724 -3434 -620 -3060
rect -4113 -3486 -991 -3485
rect -4113 -6606 -4112 -3486
rect -992 -6606 -991 -3486
rect -4113 -6607 -991 -6606
rect -2604 -7083 -2500 -6607
rect -724 -6658 -704 -3434
rect -640 -6658 -620 -3434
rect 1708 -3485 1812 -3009
rect 3588 -3060 3608 164
rect 3672 -3060 3692 164
rect 3588 -3434 3692 -3060
rect 199 -3486 3321 -3485
rect 199 -6606 200 -3486
rect 3320 -6606 3321 -3486
rect 199 -6607 3321 -6606
rect -724 -7032 -620 -6658
rect -4113 -7084 -991 -7083
rect -4113 -10204 -4112 -7084
rect -992 -10204 -991 -7084
rect -4113 -10205 -991 -10204
rect -2604 -10681 -2500 -10205
rect -724 -10256 -704 -7032
rect -640 -10256 -620 -7032
rect 1708 -7083 1812 -6607
rect 3588 -6658 3608 -3434
rect 3672 -6658 3692 -3434
rect 3588 -7032 3692 -6658
rect 199 -7084 3321 -7083
rect 199 -10204 200 -7084
rect 3320 -10204 3321 -7084
rect 199 -10205 3321 -10204
rect -724 -10630 -620 -10256
rect -4113 -10682 -991 -10681
rect -4113 -13802 -4112 -10682
rect -992 -13802 -991 -10682
rect -4113 -13803 -991 -13802
rect -2604 -14279 -2500 -13803
rect -724 -13854 -704 -10630
rect -640 -13854 -620 -10630
rect 1708 -10681 1812 -10205
rect 3588 -10256 3608 -7032
rect 3672 -10256 3692 -7032
rect 3588 -10630 3692 -10256
rect 199 -10682 3321 -10681
rect 199 -13802 200 -10682
rect 3320 -13802 3321 -10682
rect 199 -13803 3321 -13802
rect -724 -14228 -620 -13854
rect -4113 -14280 -991 -14279
rect -4113 -17400 -4112 -14280
rect -992 -17400 -991 -14280
rect -4113 -17401 -991 -17400
rect -2604 -17600 -2500 -17401
rect -724 -17452 -704 -14228
rect -640 -17452 -620 -14228
rect 1708 -14279 1812 -13803
rect 3588 -13854 3608 -10630
rect 3672 -13854 3692 -10630
rect 3588 -14228 3692 -13854
rect 199 -14280 3321 -14279
rect 199 -17400 200 -14280
rect 3320 -17400 3321 -14280
rect 199 -17401 3321 -17400
rect -724 -17600 -620 -17452
rect 1708 -17600 1812 -17401
rect 3588 -17452 3608 -14228
rect 3672 -17452 3692 -14228
rect 3588 -17600 3692 -17452
<< properties >>
string FIXED_BBOX 120 14200 3400 17480
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 16.00 l 16.00 val 524.159 carea 2.00 cperi 0.19 nx 2 ny 10 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
