magic
tech sky130A
magscale 1 2
timestamp 1717527227
<< pwell >>
rect -318 -567 318 567
<< mvnnmos >>
rect -90 109 90 309
rect -90 -309 90 -109
<< mvndiff >>
rect -148 297 -90 309
rect -148 121 -136 297
rect -102 121 -90 297
rect -148 109 -90 121
rect 90 297 148 309
rect 90 121 102 297
rect 136 121 148 297
rect 90 109 148 121
rect -148 -121 -90 -109
rect -148 -297 -136 -121
rect -102 -297 -90 -121
rect -148 -309 -90 -297
rect 90 -121 148 -109
rect 90 -297 102 -121
rect 136 -297 148 -121
rect 90 -309 148 -297
<< mvndiffc >>
rect -136 121 -102 297
rect 102 121 136 297
rect -136 -297 -102 -121
rect 102 -297 136 -121
<< mvpsubdiff >>
rect -282 519 282 531
rect -282 485 -174 519
rect 174 485 282 519
rect -282 473 282 485
rect -282 423 -224 473
rect -282 -423 -270 423
rect -236 -423 -224 423
rect 224 423 282 473
rect -282 -473 -224 -423
rect 224 -423 236 423
rect 270 -423 282 423
rect 224 -473 282 -423
rect -282 -485 282 -473
rect -282 -519 -174 -485
rect 174 -519 282 -485
rect -282 -531 282 -519
<< mvpsubdiffcont >>
rect -174 485 174 519
rect -270 -423 -236 423
rect 236 -423 270 423
rect -174 -519 174 -485
<< poly >>
rect -90 381 90 397
rect -90 347 -74 381
rect 74 347 90 381
rect -90 309 90 347
rect -90 71 90 109
rect -90 37 -74 71
rect 74 37 90 71
rect -90 21 90 37
rect -90 -37 90 -21
rect -90 -71 -74 -37
rect 74 -71 90 -37
rect -90 -109 90 -71
rect -90 -347 90 -309
rect -90 -381 -74 -347
rect 74 -381 90 -347
rect -90 -397 90 -381
<< polycont >>
rect -74 347 74 381
rect -74 37 74 71
rect -74 -71 74 -37
rect -74 -381 74 -347
<< locali >>
rect -270 485 -174 519
rect 174 485 270 519
rect -270 423 -236 485
rect 236 423 270 485
rect -90 347 -74 381
rect 74 347 90 381
rect -136 297 -102 313
rect -136 105 -102 121
rect 102 297 136 313
rect 102 105 136 121
rect -90 37 -74 71
rect 74 37 90 71
rect -90 -71 -74 -37
rect 74 -71 90 -37
rect -136 -121 -102 -105
rect -136 -313 -102 -297
rect 102 -121 136 -105
rect 102 -313 136 -297
rect -90 -381 -74 -347
rect 74 -381 90 -347
rect -270 -485 -236 -423
rect 236 -485 270 -423
rect -270 -519 -174 -485
rect 174 -519 270 -485
<< viali >>
rect -74 347 74 381
rect -136 121 -102 297
rect 102 121 136 297
rect -74 37 74 71
rect -74 -71 74 -37
rect -136 -297 -102 -121
rect 102 -297 136 -121
rect -74 -381 74 -347
<< metal1 >>
rect -86 381 86 387
rect -86 347 -74 381
rect 74 347 86 381
rect -86 341 86 347
rect -142 297 -96 309
rect -142 121 -136 297
rect -102 121 -96 297
rect -142 109 -96 121
rect 96 297 142 309
rect 96 121 102 297
rect 136 121 142 297
rect 96 109 142 121
rect -86 71 86 77
rect -86 37 -74 71
rect 74 37 86 71
rect -86 31 86 37
rect -86 -37 86 -31
rect -86 -71 -74 -37
rect 74 -71 86 -37
rect -86 -77 86 -71
rect -142 -121 -96 -109
rect -142 -297 -136 -121
rect -102 -297 -96 -121
rect -142 -309 -96 -297
rect 96 -121 142 -109
rect 96 -297 102 -121
rect 136 -297 142 -121
rect 96 -309 142 -297
rect -86 -347 86 -341
rect -86 -381 -74 -347
rect 74 -381 86 -347
rect -86 -387 86 -381
<< properties >>
string FIXED_BBOX -253 -502 253 502
string gencell sky130_fd_pr__nfet_05v0_nvt
string library sky130
string parameters w 1.0 l 0.9 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.90 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
