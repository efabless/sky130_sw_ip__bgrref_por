magic
tech sky130A
timestamp 1717527227
<< pwell >>
rect -159 -229 159 229
<< mvnmos >>
rect -40 -100 40 100
<< mvndiff >>
rect -69 94 -40 100
rect -69 -94 -63 94
rect -46 -94 -40 94
rect -69 -100 -40 -94
rect 40 94 69 100
rect 40 -94 46 94
rect 63 -94 69 94
rect 40 -100 69 -94
<< mvndiffc >>
rect -63 -94 -46 94
rect 46 -94 63 94
<< mvpsubdiff >>
rect -141 205 141 211
rect -141 188 -82 205
rect 82 188 141 205
rect -141 182 141 188
rect -141 157 -112 182
rect -141 -157 -135 157
rect -118 -157 -112 157
rect 112 157 141 182
rect -141 -182 -112 -157
rect 112 -157 118 157
rect 135 -157 141 157
rect 112 -182 141 -157
rect -141 -188 141 -182
rect -141 -205 -82 -188
rect 82 -205 141 -188
rect -141 -211 141 -205
<< mvpsubdiffcont >>
rect -82 188 82 205
rect -135 -157 -118 157
rect 118 -157 135 157
rect -82 -205 82 -188
<< poly >>
rect -40 136 40 144
rect -40 119 -32 136
rect 32 119 40 136
rect -40 100 40 119
rect -40 -119 40 -100
rect -40 -136 -32 -119
rect 32 -136 40 -119
rect -40 -144 40 -136
<< polycont >>
rect -32 119 32 136
rect -32 -136 32 -119
<< locali >>
rect -135 188 -82 205
rect 82 188 135 205
rect -135 157 -118 188
rect 118 157 135 188
rect -40 119 -32 136
rect 32 119 40 136
rect -63 94 -46 102
rect -63 -102 -46 -94
rect 46 94 63 102
rect 46 -102 63 -94
rect -40 -136 -32 -119
rect 32 -136 40 -119
rect -135 -188 -118 -157
rect 118 -188 135 -157
rect -135 -205 -82 -188
rect 82 -205 135 -188
<< viali >>
rect -32 119 32 136
rect -63 -94 -46 94
rect 46 -94 63 94
rect -32 -136 32 -119
<< metal1 >>
rect -38 136 38 139
rect -38 119 -32 136
rect 32 119 38 136
rect -38 116 38 119
rect -66 94 -43 100
rect -66 -94 -63 94
rect -46 -94 -43 94
rect -66 -100 -43 -94
rect 43 94 66 100
rect 43 -94 46 94
rect 63 -94 66 94
rect 43 -100 66 -94
rect -38 -119 38 -116
rect -38 -136 -32 -119
rect 32 -136 38 -119
rect -38 -139 38 -136
<< properties >>
string FIXED_BBOX -121 -196 121 196
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2.0 l 0.8 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
