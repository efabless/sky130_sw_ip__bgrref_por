magic
tech sky130A
magscale 1 2
timestamp 1731359787
<< pwell >>
rect -1363 -4582 1363 4582
<< psubdiff >>
rect -1327 4512 -1231 4546
rect 1231 4512 1327 4546
rect -1327 4450 -1293 4512
rect 1293 4450 1327 4512
rect -1327 -4512 -1293 -4450
rect 1293 -4512 1327 -4450
rect -1327 -4546 -1231 -4512
rect 1231 -4546 1327 -4512
<< psubdiffcont >>
rect -1231 4512 1231 4546
rect -1327 -4450 -1293 4450
rect 1293 -4450 1327 4450
rect -1231 -4546 1231 -4512
<< xpolycontact >>
rect -1197 3984 -1127 4416
rect -1197 -4416 -1127 -3984
rect -1031 3984 -961 4416
rect -1031 -4416 -961 -3984
rect -865 3984 -795 4416
rect -865 -4416 -795 -3984
rect -699 3984 -629 4416
rect -699 -4416 -629 -3984
rect -533 3984 -463 4416
rect -533 -4416 -463 -3984
rect -367 3984 -297 4416
rect -367 -4416 -297 -3984
rect -201 3984 -131 4416
rect -201 -4416 -131 -3984
rect -35 3984 35 4416
rect -35 -4416 35 -3984
rect 131 3984 201 4416
rect 131 -4416 201 -3984
rect 297 3984 367 4416
rect 297 -4416 367 -3984
rect 463 3984 533 4416
rect 463 -4416 533 -3984
rect 629 3984 699 4416
rect 629 -4416 699 -3984
rect 795 3984 865 4416
rect 795 -4416 865 -3984
rect 961 3984 1031 4416
rect 961 -4416 1031 -3984
rect 1127 3984 1197 4416
rect 1127 -4416 1197 -3984
<< xpolyres >>
rect -1197 -3984 -1127 3984
rect -1031 -3984 -961 3984
rect -865 -3984 -795 3984
rect -699 -3984 -629 3984
rect -533 -3984 -463 3984
rect -367 -3984 -297 3984
rect -201 -3984 -131 3984
rect -35 -3984 35 3984
rect 131 -3984 201 3984
rect 297 -3984 367 3984
rect 463 -3984 533 3984
rect 629 -3984 699 3984
rect 795 -3984 865 3984
rect 961 -3984 1031 3984
rect 1127 -3984 1197 3984
<< locali >>
rect -1327 4512 -1231 4546
rect 1231 4512 1327 4546
rect -1327 4450 -1293 4512
rect 1293 4450 1327 4512
rect -1327 -4512 -1293 -4450
rect 1293 -4512 1327 -4450
rect -1327 -4546 -1231 -4512
rect 1231 -4546 1327 -4512
<< viali >>
rect -1181 4001 -1143 4398
rect -1015 4001 -977 4398
rect -849 4001 -811 4398
rect -683 4001 -645 4398
rect -517 4001 -479 4398
rect -351 4001 -313 4398
rect -185 4001 -147 4398
rect -19 4001 19 4398
rect 147 4001 185 4398
rect 313 4001 351 4398
rect 479 4001 517 4398
rect 645 4001 683 4398
rect 811 4001 849 4398
rect 977 4001 1015 4398
rect 1143 4001 1181 4398
rect -1181 -4398 -1143 -4001
rect -1015 -4398 -977 -4001
rect -849 -4398 -811 -4001
rect -683 -4398 -645 -4001
rect -517 -4398 -479 -4001
rect -351 -4398 -313 -4001
rect -185 -4398 -147 -4001
rect -19 -4398 19 -4001
rect 147 -4398 185 -4001
rect 313 -4398 351 -4001
rect 479 -4398 517 -4001
rect 645 -4398 683 -4001
rect 811 -4398 849 -4001
rect 977 -4398 1015 -4001
rect 1143 -4398 1181 -4001
<< metal1 >>
rect -1187 4398 -1137 4410
rect -1187 4001 -1181 4398
rect -1143 4001 -1137 4398
rect -1187 3989 -1137 4001
rect -1021 4398 -971 4410
rect -1021 4001 -1015 4398
rect -977 4001 -971 4398
rect -1021 3989 -971 4001
rect -855 4398 -805 4410
rect -855 4001 -849 4398
rect -811 4001 -805 4398
rect -855 3989 -805 4001
rect -689 4398 -639 4410
rect -689 4001 -683 4398
rect -645 4001 -639 4398
rect -689 3989 -639 4001
rect -523 4398 -473 4410
rect -523 4001 -517 4398
rect -479 4001 -473 4398
rect -523 3989 -473 4001
rect -357 4398 -307 4410
rect -357 4001 -351 4398
rect -313 4001 -307 4398
rect -357 3989 -307 4001
rect -191 4398 -141 4410
rect -191 4001 -185 4398
rect -147 4001 -141 4398
rect -191 3989 -141 4001
rect -25 4398 25 4410
rect -25 4001 -19 4398
rect 19 4001 25 4398
rect -25 3989 25 4001
rect 141 4398 191 4410
rect 141 4001 147 4398
rect 185 4001 191 4398
rect 141 3989 191 4001
rect 307 4398 357 4410
rect 307 4001 313 4398
rect 351 4001 357 4398
rect 307 3989 357 4001
rect 473 4398 523 4410
rect 473 4001 479 4398
rect 517 4001 523 4398
rect 473 3989 523 4001
rect 639 4398 689 4410
rect 639 4001 645 4398
rect 683 4001 689 4398
rect 639 3989 689 4001
rect 805 4398 855 4410
rect 805 4001 811 4398
rect 849 4001 855 4398
rect 805 3989 855 4001
rect 971 4398 1021 4410
rect 971 4001 977 4398
rect 1015 4001 1021 4398
rect 971 3989 1021 4001
rect 1137 4398 1187 4410
rect 1137 4001 1143 4398
rect 1181 4001 1187 4398
rect 1137 3989 1187 4001
rect -1187 -4001 -1137 -3989
rect -1187 -4398 -1181 -4001
rect -1143 -4398 -1137 -4001
rect -1187 -4410 -1137 -4398
rect -1021 -4001 -971 -3989
rect -1021 -4398 -1015 -4001
rect -977 -4398 -971 -4001
rect -1021 -4410 -971 -4398
rect -855 -4001 -805 -3989
rect -855 -4398 -849 -4001
rect -811 -4398 -805 -4001
rect -855 -4410 -805 -4398
rect -689 -4001 -639 -3989
rect -689 -4398 -683 -4001
rect -645 -4398 -639 -4001
rect -689 -4410 -639 -4398
rect -523 -4001 -473 -3989
rect -523 -4398 -517 -4001
rect -479 -4398 -473 -4001
rect -523 -4410 -473 -4398
rect -357 -4001 -307 -3989
rect -357 -4398 -351 -4001
rect -313 -4398 -307 -4001
rect -357 -4410 -307 -4398
rect -191 -4001 -141 -3989
rect -191 -4398 -185 -4001
rect -147 -4398 -141 -4001
rect -191 -4410 -141 -4398
rect -25 -4001 25 -3989
rect -25 -4398 -19 -4001
rect 19 -4398 25 -4001
rect -25 -4410 25 -4398
rect 141 -4001 191 -3989
rect 141 -4398 147 -4001
rect 185 -4398 191 -4001
rect 141 -4410 191 -4398
rect 307 -4001 357 -3989
rect 307 -4398 313 -4001
rect 351 -4398 357 -4001
rect 307 -4410 357 -4398
rect 473 -4001 523 -3989
rect 473 -4398 479 -4001
rect 517 -4398 523 -4001
rect 473 -4410 523 -4398
rect 639 -4001 689 -3989
rect 639 -4398 645 -4001
rect 683 -4398 689 -4001
rect 639 -4410 689 -4398
rect 805 -4001 855 -3989
rect 805 -4398 811 -4001
rect 849 -4398 855 -4001
rect 805 -4410 855 -4398
rect 971 -4001 1021 -3989
rect 971 -4398 977 -4001
rect 1015 -4398 1021 -4001
rect 971 -4410 1021 -4398
rect 1137 -4001 1187 -3989
rect 1137 -4398 1143 -4001
rect 1181 -4398 1187 -4001
rect 1137 -4410 1187 -4398
<< properties >>
string FIXED_BBOX -1310 -4529 1310 4529
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 40 m 1 nx 15 wmin 0.350 lmin 0.50 class resistor rho 2000 val 229.646k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
