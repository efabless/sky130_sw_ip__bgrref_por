magic
tech sky130A
magscale 1 2
timestamp 1717363523
<< error_p >>
rect -77 1467 -19 1473
rect -77 1433 -65 1467
rect -77 1427 -19 1433
rect 19 1199 77 1205
rect 19 1165 31 1199
rect 19 1159 77 1165
rect 19 1091 77 1097
rect 19 1057 31 1091
rect 19 1051 77 1057
rect -77 823 -19 829
rect -77 789 -65 823
rect -77 783 -19 789
rect -77 715 -19 721
rect -77 681 -65 715
rect -77 675 -19 681
rect 19 447 77 453
rect 19 413 31 447
rect 19 407 77 413
rect 19 339 77 345
rect 19 305 31 339
rect 19 299 77 305
rect -77 71 -19 77
rect -77 37 -65 71
rect -77 31 -19 37
rect -77 -37 -19 -31
rect -77 -71 -65 -37
rect -77 -77 -19 -71
rect 19 -305 77 -299
rect 19 -339 31 -305
rect 19 -345 77 -339
rect 19 -413 77 -407
rect 19 -447 31 -413
rect 19 -453 77 -447
rect -77 -681 -19 -675
rect -77 -715 -65 -681
rect -77 -721 -19 -715
rect -77 -789 -19 -783
rect -77 -823 -65 -789
rect -77 -829 -19 -823
rect 19 -1057 77 -1051
rect 19 -1091 31 -1057
rect 19 -1097 77 -1091
rect 19 -1165 77 -1159
rect 19 -1199 31 -1165
rect 19 -1205 77 -1199
rect -77 -1433 -19 -1427
rect -77 -1467 -65 -1433
rect -77 -1473 -19 -1467
<< nwell >>
rect -263 -1605 263 1605
<< pmos >>
rect -63 1246 -33 1386
rect 33 1246 63 1386
rect -63 870 -33 1010
rect 33 870 63 1010
rect -63 494 -33 634
rect 33 494 63 634
rect -63 118 -33 258
rect 33 118 63 258
rect -63 -258 -33 -118
rect 33 -258 63 -118
rect -63 -634 -33 -494
rect 33 -634 63 -494
rect -63 -1010 -33 -870
rect 33 -1010 63 -870
rect -63 -1386 -33 -1246
rect 33 -1386 63 -1246
<< pdiff >>
rect -125 1374 -63 1386
rect -125 1258 -113 1374
rect -79 1258 -63 1374
rect -125 1246 -63 1258
rect -33 1374 33 1386
rect -33 1258 -17 1374
rect 17 1258 33 1374
rect -33 1246 33 1258
rect 63 1374 125 1386
rect 63 1258 79 1374
rect 113 1258 125 1374
rect 63 1246 125 1258
rect -125 998 -63 1010
rect -125 882 -113 998
rect -79 882 -63 998
rect -125 870 -63 882
rect -33 998 33 1010
rect -33 882 -17 998
rect 17 882 33 998
rect -33 870 33 882
rect 63 998 125 1010
rect 63 882 79 998
rect 113 882 125 998
rect 63 870 125 882
rect -125 622 -63 634
rect -125 506 -113 622
rect -79 506 -63 622
rect -125 494 -63 506
rect -33 622 33 634
rect -33 506 -17 622
rect 17 506 33 622
rect -33 494 33 506
rect 63 622 125 634
rect 63 506 79 622
rect 113 506 125 622
rect 63 494 125 506
rect -125 246 -63 258
rect -125 130 -113 246
rect -79 130 -63 246
rect -125 118 -63 130
rect -33 246 33 258
rect -33 130 -17 246
rect 17 130 33 246
rect -33 118 33 130
rect 63 246 125 258
rect 63 130 79 246
rect 113 130 125 246
rect 63 118 125 130
rect -125 -130 -63 -118
rect -125 -246 -113 -130
rect -79 -246 -63 -130
rect -125 -258 -63 -246
rect -33 -130 33 -118
rect -33 -246 -17 -130
rect 17 -246 33 -130
rect -33 -258 33 -246
rect 63 -130 125 -118
rect 63 -246 79 -130
rect 113 -246 125 -130
rect 63 -258 125 -246
rect -125 -506 -63 -494
rect -125 -622 -113 -506
rect -79 -622 -63 -506
rect -125 -634 -63 -622
rect -33 -506 33 -494
rect -33 -622 -17 -506
rect 17 -622 33 -506
rect -33 -634 33 -622
rect 63 -506 125 -494
rect 63 -622 79 -506
rect 113 -622 125 -506
rect 63 -634 125 -622
rect -125 -882 -63 -870
rect -125 -998 -113 -882
rect -79 -998 -63 -882
rect -125 -1010 -63 -998
rect -33 -882 33 -870
rect -33 -998 -17 -882
rect 17 -998 33 -882
rect -33 -1010 33 -998
rect 63 -882 125 -870
rect 63 -998 79 -882
rect 113 -998 125 -882
rect 63 -1010 125 -998
rect -125 -1258 -63 -1246
rect -125 -1374 -113 -1258
rect -79 -1374 -63 -1258
rect -125 -1386 -63 -1374
rect -33 -1258 33 -1246
rect -33 -1374 -17 -1258
rect 17 -1374 33 -1258
rect -33 -1386 33 -1374
rect 63 -1258 125 -1246
rect 63 -1374 79 -1258
rect 113 -1374 125 -1258
rect 63 -1386 125 -1374
<< pdiffc >>
rect -113 1258 -79 1374
rect -17 1258 17 1374
rect 79 1258 113 1374
rect -113 882 -79 998
rect -17 882 17 998
rect 79 882 113 998
rect -113 506 -79 622
rect -17 506 17 622
rect 79 506 113 622
rect -113 130 -79 246
rect -17 130 17 246
rect 79 130 113 246
rect -113 -246 -79 -130
rect -17 -246 17 -130
rect 79 -246 113 -130
rect -113 -622 -79 -506
rect -17 -622 17 -506
rect 79 -622 113 -506
rect -113 -998 -79 -882
rect -17 -998 17 -882
rect 79 -998 113 -882
rect -113 -1374 -79 -1258
rect -17 -1374 17 -1258
rect 79 -1374 113 -1258
<< nsubdiff >>
rect -227 1535 -131 1569
rect 131 1535 227 1569
rect -227 1473 -193 1535
rect 193 1473 227 1535
rect -227 -1535 -193 -1473
rect 193 -1535 227 -1473
rect -227 -1569 -131 -1535
rect 131 -1569 227 -1535
<< nsubdiffcont >>
rect -131 1535 131 1569
rect -227 -1473 -193 1473
rect 193 -1473 227 1473
rect -131 -1569 131 -1535
<< poly >>
rect -81 1467 -15 1483
rect -81 1433 -65 1467
rect -31 1433 -15 1467
rect -81 1417 -15 1433
rect -63 1386 -33 1417
rect 33 1386 63 1412
rect -63 1220 -33 1246
rect 33 1215 63 1246
rect 15 1199 81 1215
rect 15 1165 31 1199
rect 65 1165 81 1199
rect 15 1149 81 1165
rect 15 1091 81 1107
rect 15 1057 31 1091
rect 65 1057 81 1091
rect 15 1041 81 1057
rect -63 1010 -33 1036
rect 33 1010 63 1041
rect -63 839 -33 870
rect 33 844 63 870
rect -81 823 -15 839
rect -81 789 -65 823
rect -31 789 -15 823
rect -81 773 -15 789
rect -81 715 -15 731
rect -81 681 -65 715
rect -31 681 -15 715
rect -81 665 -15 681
rect -63 634 -33 665
rect 33 634 63 660
rect -63 468 -33 494
rect 33 463 63 494
rect 15 447 81 463
rect 15 413 31 447
rect 65 413 81 447
rect 15 397 81 413
rect 15 339 81 355
rect 15 305 31 339
rect 65 305 81 339
rect 15 289 81 305
rect -63 258 -33 284
rect 33 258 63 289
rect -63 87 -33 118
rect 33 92 63 118
rect -81 71 -15 87
rect -81 37 -65 71
rect -31 37 -15 71
rect -81 21 -15 37
rect -81 -37 -15 -21
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect -81 -87 -15 -71
rect -63 -118 -33 -87
rect 33 -118 63 -92
rect -63 -284 -33 -258
rect 33 -289 63 -258
rect 15 -305 81 -289
rect 15 -339 31 -305
rect 65 -339 81 -305
rect 15 -355 81 -339
rect 15 -413 81 -397
rect 15 -447 31 -413
rect 65 -447 81 -413
rect 15 -463 81 -447
rect -63 -494 -33 -468
rect 33 -494 63 -463
rect -63 -665 -33 -634
rect 33 -660 63 -634
rect -81 -681 -15 -665
rect -81 -715 -65 -681
rect -31 -715 -15 -681
rect -81 -731 -15 -715
rect -81 -789 -15 -773
rect -81 -823 -65 -789
rect -31 -823 -15 -789
rect -81 -839 -15 -823
rect -63 -870 -33 -839
rect 33 -870 63 -844
rect -63 -1036 -33 -1010
rect 33 -1041 63 -1010
rect 15 -1057 81 -1041
rect 15 -1091 31 -1057
rect 65 -1091 81 -1057
rect 15 -1107 81 -1091
rect 15 -1165 81 -1149
rect 15 -1199 31 -1165
rect 65 -1199 81 -1165
rect 15 -1215 81 -1199
rect -63 -1246 -33 -1220
rect 33 -1246 63 -1215
rect -63 -1417 -33 -1386
rect 33 -1412 63 -1386
rect -81 -1433 -15 -1417
rect -81 -1467 -65 -1433
rect -31 -1467 -15 -1433
rect -81 -1483 -15 -1467
<< polycont >>
rect -65 1433 -31 1467
rect 31 1165 65 1199
rect 31 1057 65 1091
rect -65 789 -31 823
rect -65 681 -31 715
rect 31 413 65 447
rect 31 305 65 339
rect -65 37 -31 71
rect -65 -71 -31 -37
rect 31 -339 65 -305
rect 31 -447 65 -413
rect -65 -715 -31 -681
rect -65 -823 -31 -789
rect 31 -1091 65 -1057
rect 31 -1199 65 -1165
rect -65 -1467 -31 -1433
<< locali >>
rect -227 1535 -131 1569
rect 131 1535 227 1569
rect -227 1473 -193 1535
rect 193 1473 227 1535
rect -81 1433 -65 1467
rect -31 1433 -15 1467
rect -113 1374 -79 1390
rect -113 1242 -79 1258
rect -17 1374 17 1390
rect -17 1242 17 1258
rect 79 1374 113 1390
rect 79 1242 113 1258
rect 15 1165 31 1199
rect 65 1165 81 1199
rect 15 1057 31 1091
rect 65 1057 81 1091
rect -113 998 -79 1014
rect -113 866 -79 882
rect -17 998 17 1014
rect -17 866 17 882
rect 79 998 113 1014
rect 79 866 113 882
rect -81 789 -65 823
rect -31 789 -15 823
rect -81 681 -65 715
rect -31 681 -15 715
rect -113 622 -79 638
rect -113 490 -79 506
rect -17 622 17 638
rect -17 490 17 506
rect 79 622 113 638
rect 79 490 113 506
rect 15 413 31 447
rect 65 413 81 447
rect 15 305 31 339
rect 65 305 81 339
rect -113 246 -79 262
rect -113 114 -79 130
rect -17 246 17 262
rect -17 114 17 130
rect 79 246 113 262
rect 79 114 113 130
rect -81 37 -65 71
rect -31 37 -15 71
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect -113 -130 -79 -114
rect -113 -262 -79 -246
rect -17 -130 17 -114
rect -17 -262 17 -246
rect 79 -130 113 -114
rect 79 -262 113 -246
rect 15 -339 31 -305
rect 65 -339 81 -305
rect 15 -447 31 -413
rect 65 -447 81 -413
rect -113 -506 -79 -490
rect -113 -638 -79 -622
rect -17 -506 17 -490
rect -17 -638 17 -622
rect 79 -506 113 -490
rect 79 -638 113 -622
rect -81 -715 -65 -681
rect -31 -715 -15 -681
rect -81 -823 -65 -789
rect -31 -823 -15 -789
rect -113 -882 -79 -866
rect -113 -1014 -79 -998
rect -17 -882 17 -866
rect -17 -1014 17 -998
rect 79 -882 113 -866
rect 79 -1014 113 -998
rect 15 -1091 31 -1057
rect 65 -1091 81 -1057
rect 15 -1199 31 -1165
rect 65 -1199 81 -1165
rect -113 -1258 -79 -1242
rect -113 -1390 -79 -1374
rect -17 -1258 17 -1242
rect -17 -1390 17 -1374
rect 79 -1258 113 -1242
rect 79 -1390 113 -1374
rect -81 -1467 -65 -1433
rect -31 -1467 -15 -1433
rect -227 -1535 -193 -1473
rect 193 -1535 227 -1473
rect -227 -1569 -131 -1535
rect 131 -1569 227 -1535
<< viali >>
rect -65 1433 -31 1467
rect -113 1258 -79 1374
rect -17 1258 17 1374
rect 79 1258 113 1374
rect 31 1165 65 1199
rect 31 1057 65 1091
rect -113 882 -79 998
rect -17 882 17 998
rect 79 882 113 998
rect -65 789 -31 823
rect -65 681 -31 715
rect -113 506 -79 622
rect -17 506 17 622
rect 79 506 113 622
rect 31 413 65 447
rect 31 305 65 339
rect -113 130 -79 246
rect -17 130 17 246
rect 79 130 113 246
rect -65 37 -31 71
rect -65 -71 -31 -37
rect -113 -246 -79 -130
rect -17 -246 17 -130
rect 79 -246 113 -130
rect 31 -339 65 -305
rect 31 -447 65 -413
rect -113 -622 -79 -506
rect -17 -622 17 -506
rect 79 -622 113 -506
rect -65 -715 -31 -681
rect -65 -823 -31 -789
rect -113 -998 -79 -882
rect -17 -998 17 -882
rect 79 -998 113 -882
rect 31 -1091 65 -1057
rect 31 -1199 65 -1165
rect -113 -1374 -79 -1258
rect -17 -1374 17 -1258
rect 79 -1374 113 -1258
rect -65 -1467 -31 -1433
<< metal1 >>
rect -77 1467 -19 1473
rect -77 1433 -65 1467
rect -31 1433 -19 1467
rect -77 1427 -19 1433
rect -119 1374 -73 1386
rect -119 1258 -113 1374
rect -79 1258 -73 1374
rect -119 1246 -73 1258
rect -23 1374 23 1386
rect -23 1258 -17 1374
rect 17 1258 23 1374
rect -23 1246 23 1258
rect 73 1374 119 1386
rect 73 1258 79 1374
rect 113 1258 119 1374
rect 73 1246 119 1258
rect 19 1199 77 1205
rect 19 1165 31 1199
rect 65 1165 77 1199
rect 19 1159 77 1165
rect 19 1091 77 1097
rect 19 1057 31 1091
rect 65 1057 77 1091
rect 19 1051 77 1057
rect -119 998 -73 1010
rect -119 882 -113 998
rect -79 882 -73 998
rect -119 870 -73 882
rect -23 998 23 1010
rect -23 882 -17 998
rect 17 882 23 998
rect -23 870 23 882
rect 73 998 119 1010
rect 73 882 79 998
rect 113 882 119 998
rect 73 870 119 882
rect -77 823 -19 829
rect -77 789 -65 823
rect -31 789 -19 823
rect -77 783 -19 789
rect -77 715 -19 721
rect -77 681 -65 715
rect -31 681 -19 715
rect -77 675 -19 681
rect -119 622 -73 634
rect -119 506 -113 622
rect -79 506 -73 622
rect -119 494 -73 506
rect -23 622 23 634
rect -23 506 -17 622
rect 17 506 23 622
rect -23 494 23 506
rect 73 622 119 634
rect 73 506 79 622
rect 113 506 119 622
rect 73 494 119 506
rect 19 447 77 453
rect 19 413 31 447
rect 65 413 77 447
rect 19 407 77 413
rect 19 339 77 345
rect 19 305 31 339
rect 65 305 77 339
rect 19 299 77 305
rect -119 246 -73 258
rect -119 130 -113 246
rect -79 130 -73 246
rect -119 118 -73 130
rect -23 246 23 258
rect -23 130 -17 246
rect 17 130 23 246
rect -23 118 23 130
rect 73 246 119 258
rect 73 130 79 246
rect 113 130 119 246
rect 73 118 119 130
rect -77 71 -19 77
rect -77 37 -65 71
rect -31 37 -19 71
rect -77 31 -19 37
rect -77 -37 -19 -31
rect -77 -71 -65 -37
rect -31 -71 -19 -37
rect -77 -77 -19 -71
rect -119 -130 -73 -118
rect -119 -246 -113 -130
rect -79 -246 -73 -130
rect -119 -258 -73 -246
rect -23 -130 23 -118
rect -23 -246 -17 -130
rect 17 -246 23 -130
rect -23 -258 23 -246
rect 73 -130 119 -118
rect 73 -246 79 -130
rect 113 -246 119 -130
rect 73 -258 119 -246
rect 19 -305 77 -299
rect 19 -339 31 -305
rect 65 -339 77 -305
rect 19 -345 77 -339
rect 19 -413 77 -407
rect 19 -447 31 -413
rect 65 -447 77 -413
rect 19 -453 77 -447
rect -119 -506 -73 -494
rect -119 -622 -113 -506
rect -79 -622 -73 -506
rect -119 -634 -73 -622
rect -23 -506 23 -494
rect -23 -622 -17 -506
rect 17 -622 23 -506
rect -23 -634 23 -622
rect 73 -506 119 -494
rect 73 -622 79 -506
rect 113 -622 119 -506
rect 73 -634 119 -622
rect -77 -681 -19 -675
rect -77 -715 -65 -681
rect -31 -715 -19 -681
rect -77 -721 -19 -715
rect -77 -789 -19 -783
rect -77 -823 -65 -789
rect -31 -823 -19 -789
rect -77 -829 -19 -823
rect -119 -882 -73 -870
rect -119 -998 -113 -882
rect -79 -998 -73 -882
rect -119 -1010 -73 -998
rect -23 -882 23 -870
rect -23 -998 -17 -882
rect 17 -998 23 -882
rect -23 -1010 23 -998
rect 73 -882 119 -870
rect 73 -998 79 -882
rect 113 -998 119 -882
rect 73 -1010 119 -998
rect 19 -1057 77 -1051
rect 19 -1091 31 -1057
rect 65 -1091 77 -1057
rect 19 -1097 77 -1091
rect 19 -1165 77 -1159
rect 19 -1199 31 -1165
rect 65 -1199 77 -1165
rect 19 -1205 77 -1199
rect -119 -1258 -73 -1246
rect -119 -1374 -113 -1258
rect -79 -1374 -73 -1258
rect -119 -1386 -73 -1374
rect -23 -1258 23 -1246
rect -23 -1374 -17 -1258
rect 17 -1374 23 -1258
rect -23 -1386 23 -1374
rect 73 -1258 119 -1246
rect 73 -1374 79 -1258
rect 113 -1374 119 -1258
rect 73 -1386 119 -1374
rect -77 -1433 -19 -1427
rect -77 -1467 -65 -1433
rect -31 -1467 -19 -1433
rect -77 -1473 -19 -1467
<< properties >>
string FIXED_BBOX -210 -1552 210 1552
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.7 l 0.15 m 8 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
