** sch_path: /home/tim/gits/cheetah_v4_analog/dependencies/sky130_sw_ip__por/xschem/sky130_sw_ip__por.sch
.subckt sky130_sw_ip__por por avss avdd dvdd porb dvss porb_h[1] porb_h[0]
*.PININFO avdd:B por:O avss:B dvdd:B porb:O porb_h[1:0]:O dvss:B
x1 Vinn Vinp RST avss net1 dvdd vo net6 comparator_final
XR1 avss Vinn avss sky130_fd_pr__res_xhigh_po_0p35 L=1000 mult=1 m=1
XR10 Vinn Vinp avss sky130_fd_pr__res_xhigh_po_0p35 L=72 mult=1 m=1
XR12 Vinp net3 avss sky130_fd_pr__res_xhigh_po_0p35 L=600 mult=1 m=1
x2 RST por dvdd dvss net2 porb porb_h[1] porb_h[0] net6 delayPulse_final
XM2 avdd avdd net4 avss sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 nf=1 m=1
Vrbranch Vproc net3 0
.save i(vrbranch)
Vcomp avdd net1 0
.save i(vcomp)
Vpulse avdd net2 0
.save i(vpulse)
XM1 net4 avdd Vproc avss sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 nf=1 m=1
XR2 net5 Vinp avss sky130_fd_pr__res_xhigh_po_0p35 L=72 mult=1 m=1
XM3 net5 vo Vinn avss sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 nf=1 m=1
.ends

* expanding   symbol:  comparator_final.sym # of pins=8
** sym_path: /home/tim/gits/cheetah_v4_analog/dependencies/sky130_sw_ip__por/xschem/comparator_final.sym
** sch_path: /home/tim/gits/cheetah_v4_analog/dependencies/sky130_sw_ip__por/xschem/comparator_final.sch
.subckt comparator_final Vinn Vinp RST VSS AVDD DVDD vo ibn180n
*.PININFO AVDD:I RST:O VSS:I Vinn:I Vinp:I DVDD:I vo:O ibn180n:O
XM1 VS vbn VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XM3 vbp vbp AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM2 vt vbp AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM7 vo vt AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM6 vo vbn VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XM14 vo1 vo VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM15 vo1 vo net1 net1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM12 net4 vo1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM13 net4 vo1 DVDD DVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM16 RST net4 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM17 RST net4 DVDD DVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM4 vbp AVDD net3 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM8 vt AVDD net2 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM19 net1 net1 AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM23 net5 net5 AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=1 nf=1 m=1
XM24 vbn net5 AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=1 nf=1 m=1
XR12 VSS net6 VSS sky130_fd_pr__res_xhigh_po_0p35 L=28 mult=1 m=1
XM25 vbn vbn VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM26 net5 vbn net6 VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XM28 net7 vbn VSS VSS sky130_fd_pr__nfet_01v8 L=0.3 W=4 nf=1 m=1
XM18 net2 Vinn VS VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 m=7
XM10 net3 Vinp VS VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 m=2
XM5 net8 net8 AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=1 nf=1 m=1
XM11 net9 net9 net8 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=1 nf=1 m=1
XM20 net7 net7 net9 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=1 nf=1 m=1
XM21 net5 net7 vbn VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM9 net10 vbn VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=1
Vbn180n ibn180n net10 0
.save i(vbn180n)
XM22 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 m=1
.ends


* expanding   symbol:  delayPulse_final.sym # of pins=8
** sym_path: /home/tim/gits/cheetah_v4_analog/dependencies/sky130_sw_ip__por/xschem/delayPulse_final.sym
** sch_path: /home/tim/gits/cheetah_v4_analog/dependencies/sky130_sw_ip__por/xschem/delayPulse_final.sch
.subckt delayPulse_final din por VCCL VSS VCCH porb porb_h[1] porb_h[0] ibn180n
*.PININFO VCCL:I VSS:I din:I por:O VCCH:I porb:O porb_h[1:0]:O ibn180n:I
x1 Td_L Td_Sd VSS VSS VCCL VCCL outxor sky130_fd_sc_ls__xor2_1
x3 porbPre porbhPre VCCL VSS VCCH levelShifter
XM2 net1 din VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 m=2
XM3 Td_S net1 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 m=2
XM5 VT2 net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=2 m=1
XM7 net1 din VSS VSS sky130_fd_pr__nfet_01v8 L=0.3 W=0.5 nf=1 m=2
XM8 Td_S net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.3 W=0.5 nf=1 m=2
XM10 VT2 net1 net10 VCCL sky130_fd_pr__pfet_01v8 L=0.3 W=2 nf=2 m=1
XM13 net4 VT3 VSS VSS sky130_fd_pr__nfet_01v8 L=0.3 W=0.5 nf=1 m=2
XM14 net4 VT3 net5 net5 sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 m=2
x4 net2 VSS VCCL TieH_1p8
XM11 vbn1 net8 net6 VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=2 nf=1 m=1
XM17 vbp1 vbn1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=2 nf=1 m=1
XM18 net6 net7 VCCH VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=2 nf=1 m=1
XM19 vbn1 vbn1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=2 nf=1 m=7
XM24 net8 net8 net7 VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=2 nf=1 m=1
XM25 net7 net7 VCCH VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=16 nf=8 m=1
XM26 VSS VSS net9 VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XM6 VT3 VT2 net3 VSS sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=2 m=1
XM12 VT3 VT2 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.3 W=2 nf=2 m=1
XM1 vbp1 vbp1 vbp1 VCCL sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=2 m=1
XM15 vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=2 m=7
XM16 net10 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=2 m=1
XM20 net10 vbp1 net10 VCCL sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=2 m=1
XM21 net3 vbn1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=2 nf=1 m=4
XM22 net5 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=2 m=4
XM23 net5 vbp1 net5 VCCL sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=2 m=1
XM27 net11 net4 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=1
XM29 net11 net4 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=1
XM30 Td_L net11 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=2
XM31 Td_L net11 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=2
XM32 net12 Td_S VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=1
XM33 net12 Td_S VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=1
XM34 net13 net12 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=1
XM35 net13 net12 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=1
XM36 Td_Sd net14 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=2
XM38 net14 net13 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=1
XM39 net14 net13 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=1
x6 outxor VSS VSS VCCL VCCL rstn sky130_fd_sc_ls__buf_8
XC4 VSS net13 sky130_fd_pr__cap_mim_m3_2 W=10 L=10 m=1
XC7 VSS VT2 sky130_fd_pr__cap_mim_m3_2 W=16 L=16 m=20
XC2 VCCL VT3 sky130_fd_pr__cap_mim_m3_2 W=16 L=16 m=20
XC8 VCCL net12 sky130_fd_pr__cap_mim_m3_2 W=10 L=10 m=1
XC9 VCCL net14 sky130_fd_pr__cap_mim_m3_2 W=10 L=10 m=1
XM40 Td_Sd net14 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=2
x5 rstn net2 Td_Sd VSS VSS VCCL VCCL porbPre sky130_fd_sc_ls__dfrtn_1
x2 Td_Sd net2 Td_Lb VSS VSS VCCL VCCL porPre sky130_fd_sc_ls__dfrtp_1
XM4 Td_Lb Td_L VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=2
XM9 Td_Lb Td_L VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=2
XC1 VSS vbn1 sky130_fd_pr__cap_mim_m3_2 W=16 L=16 m=1
XC5 VCCH net7 sky130_fd_pr__cap_mim_m3_2 W=16 L=16 m=1
XC6 VCCL vbp1 sky130_fd_pr__cap_mim_m3_2 W=16 L=16 m=1
XC3 VCCH net8 sky130_fd_pr__cap_mim_m3_2 W=8 L=8 m=1
XM28 net15 porPre VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=1
XM37 net15 porPre VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=1
XM41 net16 net15 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=2
XM42 net16 net15 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=2
XM43 net17 net16 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=8
XM44 net17 net16 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=8
XM45 por net17 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=16
XM46 por net17 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=16
XM47 net18 porbPre VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=1
XM48 net18 porbPre VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=1
XM49 net19 net18 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=2
XM50 net19 net18 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=2
XM51 net20 net19 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=8
XM52 net20 net19 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=8
XM53 porb net20 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=16
XM54 porb net20 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=16
XM59 net21 porbhPre VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM60 net21 porbhPre VCCH VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=2 m=1
x7 VSS VSS VCCL VCCL sky130_fd_sc_ls__decap_4
XC10 net8 VCCH sky130_fd_pr__cap_mim_m3_1 W=8 L=8 m=1
XC11 net7 VCCH sky130_fd_pr__cap_mim_m3_1 W=16 L=16 m=1
XC12 vbp1 VCCL sky130_fd_pr__cap_mim_m3_1 W=16 L=16 m=1
XC13 vbn1 VSS sky130_fd_pr__cap_mim_m3_1 W=16 L=16 m=1
XC14 VT2 VSS sky130_fd_pr__cap_mim_m3_1 W=16 L=16 m=20
XC15 VT3 VCCL sky130_fd_pr__cap_mim_m3_1 W=16 L=16 m=20
XC16 net12 VCCL sky130_fd_pr__cap_mim_m3_1 W=10 L=10 m=1
XC17 net13 VSS sky130_fd_pr__cap_mim_m3_1 W=10 L=10 m=1
XC18 net14 VCCL sky130_fd_pr__cap_mim_m3_1 W=10 L=10 m=1
XR1 net23 net9 VSS sky130_fd_pr__res_xhigh_po_0p69 L=240 mult=1 m=1
XR7 VSS net23 VSS sky130_fd_pr__res_xhigh_po_0p69 L=240 mult=1 m=1
XM55 net22 net21 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM56 net22 net21 VCCH VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=2 m=1
XM57 por_h net22 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM58 por_h net22 VCCH VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=2 m=1
x10 por_h VSS VSS VCCH VCCH porb_h[0] sky130_fd_sc_hvl__inv_16
x8 por_h VSS VSS VCCH VCCH porb_h[1] sky130_fd_sc_hvl__inv_16
Vvgbias net8 ibn180n 0
.save i(vvgbias)
.ends


* expanding   symbol:  levelShifter.sym # of pins=5
** sym_path: /home/tim/gits/cheetah_v4_analog/dependencies/sky130_sw_ip__por/xschem/levelShifter.sym
** sch_path: /home/tim/gits/cheetah_v4_analog/dependencies/sky130_sw_ip__por/xschem/levelShifter.sch
.subckt levelShifter ain aout VCCL VSS VCCH
*.PININFO VCCL:I VSS:I ain:I aout:O VCCH:I
XM12 net1 S1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3.6 nf=1 m=1
XM13 aob net1 VCCH VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5.8 nf=2 m=1
XM6 S1 ain VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=1
XM1 S1 ain VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=1
XM2 net1 aob VCCH VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5.8 nf=2 m=1
XM3 aob S1B VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3.6 nf=1 m=1
XM4 S1B S1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=1
XM5 S1B S1 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=1
XM7 aout aob VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.8 nf=1 m=1
XM8 aout aob VCCH VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5.8 nf=2 m=1
XC1 VCCH aob sky130_fd_pr__cap_mim_m3_1 W=2 L=2 m=1
.ends


* expanding   symbol:  TieH_1p8.sym # of pins=3
** sym_path: /home/tim/gits/cheetah_v4_analog/dependencies/sky130_sw_ip__por/xschem/TieH_1p8.sym
** sch_path: /home/tim/gits/cheetah_v4_analog/dependencies/sky130_sw_ip__por/xschem/TieH_1p8.sch
.subckt TieH_1p8 TieH VSS VCC
*.PININFO VCC:I VSS:I TieH:B
XM4 net1 net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=1
XM5 TieH net1 VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=2 m=1
.ends

.end
