magic
tech sky130A
magscale 1 2
timestamp 1717438235
<< metal4 >>
rect -8396 8839 -4498 8880
rect -8396 5561 -4754 8839
rect -4518 5561 -4498 8839
rect -8396 5520 -4498 5561
rect -4098 8839 -200 8880
rect -4098 5561 -456 8839
rect -220 5561 -200 8839
rect -4098 5520 -200 5561
rect 200 8839 4098 8880
rect 200 5561 3842 8839
rect 4078 5561 4098 8839
rect 200 5520 4098 5561
rect 4498 8839 8396 8880
rect 4498 5561 8140 8839
rect 8376 5561 8396 8839
rect 4498 5520 8396 5561
rect -8396 5239 -4498 5280
rect -8396 1961 -4754 5239
rect -4518 1961 -4498 5239
rect -8396 1920 -4498 1961
rect -4098 5239 -200 5280
rect -4098 1961 -456 5239
rect -220 1961 -200 5239
rect -4098 1920 -200 1961
rect 200 5239 4098 5280
rect 200 1961 3842 5239
rect 4078 1961 4098 5239
rect 200 1920 4098 1961
rect 4498 5239 8396 5280
rect 4498 1961 8140 5239
rect 8376 1961 8396 5239
rect 4498 1920 8396 1961
rect -8396 1639 -4498 1680
rect -8396 -1639 -4754 1639
rect -4518 -1639 -4498 1639
rect -8396 -1680 -4498 -1639
rect -4098 1639 -200 1680
rect -4098 -1639 -456 1639
rect -220 -1639 -200 1639
rect -4098 -1680 -200 -1639
rect 200 1639 4098 1680
rect 200 -1639 3842 1639
rect 4078 -1639 4098 1639
rect 200 -1680 4098 -1639
rect 4498 1639 8396 1680
rect 4498 -1639 8140 1639
rect 8376 -1639 8396 1639
rect 4498 -1680 8396 -1639
rect -8396 -1961 -4498 -1920
rect -8396 -5239 -4754 -1961
rect -4518 -5239 -4498 -1961
rect -8396 -5280 -4498 -5239
rect -4098 -1961 -200 -1920
rect -4098 -5239 -456 -1961
rect -220 -5239 -200 -1961
rect -4098 -5280 -200 -5239
rect 200 -1961 4098 -1920
rect 200 -5239 3842 -1961
rect 4078 -5239 4098 -1961
rect 200 -5280 4098 -5239
rect 4498 -1961 8396 -1920
rect 4498 -5239 8140 -1961
rect 8376 -5239 8396 -1961
rect 4498 -5280 8396 -5239
rect -8396 -5561 -4498 -5520
rect -8396 -8839 -4754 -5561
rect -4518 -8839 -4498 -5561
rect -8396 -8880 -4498 -8839
rect -4098 -5561 -200 -5520
rect -4098 -8839 -456 -5561
rect -220 -8839 -200 -5561
rect -4098 -8880 -200 -8839
rect 200 -5561 4098 -5520
rect 200 -8839 3842 -5561
rect 4078 -8839 4098 -5561
rect 200 -8880 4098 -8839
rect 4498 -5561 8396 -5520
rect 4498 -8839 8140 -5561
rect 8376 -8839 8396 -5561
rect 4498 -8880 8396 -8839
<< via4 >>
rect -4754 5561 -4518 8839
rect -456 5561 -220 8839
rect 3842 5561 4078 8839
rect 8140 5561 8376 8839
rect -4754 1961 -4518 5239
rect -456 1961 -220 5239
rect 3842 1961 4078 5239
rect 8140 1961 8376 5239
rect -4754 -1639 -4518 1639
rect -456 -1639 -220 1639
rect 3842 -1639 4078 1639
rect 8140 -1639 8376 1639
rect -4754 -5239 -4518 -1961
rect -456 -5239 -220 -1961
rect 3842 -5239 4078 -1961
rect 8140 -5239 8376 -1961
rect -4754 -8839 -4518 -5561
rect -456 -8839 -220 -5561
rect 3842 -8839 4078 -5561
rect 8140 -8839 8376 -5561
<< mimcap2 >>
rect -8316 8760 -5116 8800
rect -8316 5640 -8276 8760
rect -5156 5640 -5116 8760
rect -8316 5600 -5116 5640
rect -4018 8760 -818 8800
rect -4018 5640 -3978 8760
rect -858 5640 -818 8760
rect -4018 5600 -818 5640
rect 280 8760 3480 8800
rect 280 5640 320 8760
rect 3440 5640 3480 8760
rect 280 5600 3480 5640
rect 4578 8760 7778 8800
rect 4578 5640 4618 8760
rect 7738 5640 7778 8760
rect 4578 5600 7778 5640
rect -8316 5160 -5116 5200
rect -8316 2040 -8276 5160
rect -5156 2040 -5116 5160
rect -8316 2000 -5116 2040
rect -4018 5160 -818 5200
rect -4018 2040 -3978 5160
rect -858 2040 -818 5160
rect -4018 2000 -818 2040
rect 280 5160 3480 5200
rect 280 2040 320 5160
rect 3440 2040 3480 5160
rect 280 2000 3480 2040
rect 4578 5160 7778 5200
rect 4578 2040 4618 5160
rect 7738 2040 7778 5160
rect 4578 2000 7778 2040
rect -8316 1560 -5116 1600
rect -8316 -1560 -8276 1560
rect -5156 -1560 -5116 1560
rect -8316 -1600 -5116 -1560
rect -4018 1560 -818 1600
rect -4018 -1560 -3978 1560
rect -858 -1560 -818 1560
rect -4018 -1600 -818 -1560
rect 280 1560 3480 1600
rect 280 -1560 320 1560
rect 3440 -1560 3480 1560
rect 280 -1600 3480 -1560
rect 4578 1560 7778 1600
rect 4578 -1560 4618 1560
rect 7738 -1560 7778 1560
rect 4578 -1600 7778 -1560
rect -8316 -2040 -5116 -2000
rect -8316 -5160 -8276 -2040
rect -5156 -5160 -5116 -2040
rect -8316 -5200 -5116 -5160
rect -4018 -2040 -818 -2000
rect -4018 -5160 -3978 -2040
rect -858 -5160 -818 -2040
rect -4018 -5200 -818 -5160
rect 280 -2040 3480 -2000
rect 280 -5160 320 -2040
rect 3440 -5160 3480 -2040
rect 280 -5200 3480 -5160
rect 4578 -2040 7778 -2000
rect 4578 -5160 4618 -2040
rect 7738 -5160 7778 -2040
rect 4578 -5200 7778 -5160
rect -8316 -5640 -5116 -5600
rect -8316 -8760 -8276 -5640
rect -5156 -8760 -5116 -5640
rect -8316 -8800 -5116 -8760
rect -4018 -5640 -818 -5600
rect -4018 -8760 -3978 -5640
rect -858 -8760 -818 -5640
rect -4018 -8800 -818 -8760
rect 280 -5640 3480 -5600
rect 280 -8760 320 -5640
rect 3440 -8760 3480 -5640
rect 280 -8800 3480 -8760
rect 4578 -5640 7778 -5600
rect 4578 -8760 4618 -5640
rect 7738 -8760 7778 -5640
rect 4578 -8800 7778 -8760
<< mimcap2contact >>
rect -8276 5640 -5156 8760
rect -3978 5640 -858 8760
rect 320 5640 3440 8760
rect 4618 5640 7738 8760
rect -8276 2040 -5156 5160
rect -3978 2040 -858 5160
rect 320 2040 3440 5160
rect 4618 2040 7738 5160
rect -8276 -1560 -5156 1560
rect -3978 -1560 -858 1560
rect 320 -1560 3440 1560
rect 4618 -1560 7738 1560
rect -8276 -5160 -5156 -2040
rect -3978 -5160 -858 -2040
rect 320 -5160 3440 -2040
rect 4618 -5160 7738 -2040
rect -8276 -8760 -5156 -5640
rect -3978 -8760 -858 -5640
rect 320 -8760 3440 -5640
rect 4618 -8760 7738 -5640
<< metal5 >>
rect -6876 8784 -6556 9000
rect -4796 8839 -4476 9000
rect -8300 8760 -5132 8784
rect -8300 5640 -8276 8760
rect -5156 5640 -5132 8760
rect -8300 5616 -5132 5640
rect -6876 5184 -6556 5616
rect -4796 5561 -4754 8839
rect -4518 5561 -4476 8839
rect -2578 8784 -2258 9000
rect -498 8839 -178 9000
rect -4002 8760 -834 8784
rect -4002 5640 -3978 8760
rect -858 5640 -834 8760
rect -4002 5616 -834 5640
rect -4796 5239 -4476 5561
rect -8300 5160 -5132 5184
rect -8300 2040 -8276 5160
rect -5156 2040 -5132 5160
rect -8300 2016 -5132 2040
rect -6876 1584 -6556 2016
rect -4796 1961 -4754 5239
rect -4518 1961 -4476 5239
rect -2578 5184 -2258 5616
rect -498 5561 -456 8839
rect -220 5561 -178 8839
rect 1720 8784 2040 9000
rect 3800 8839 4120 9000
rect 296 8760 3464 8784
rect 296 5640 320 8760
rect 3440 5640 3464 8760
rect 296 5616 3464 5640
rect -498 5239 -178 5561
rect -4002 5160 -834 5184
rect -4002 2040 -3978 5160
rect -858 2040 -834 5160
rect -4002 2016 -834 2040
rect -4796 1639 -4476 1961
rect -8300 1560 -5132 1584
rect -8300 -1560 -8276 1560
rect -5156 -1560 -5132 1560
rect -8300 -1584 -5132 -1560
rect -6876 -2016 -6556 -1584
rect -4796 -1639 -4754 1639
rect -4518 -1639 -4476 1639
rect -2578 1584 -2258 2016
rect -498 1961 -456 5239
rect -220 1961 -178 5239
rect 1720 5184 2040 5616
rect 3800 5561 3842 8839
rect 4078 5561 4120 8839
rect 6018 8784 6338 9000
rect 8098 8839 8418 9000
rect 4594 8760 7762 8784
rect 4594 5640 4618 8760
rect 7738 5640 7762 8760
rect 4594 5616 7762 5640
rect 3800 5239 4120 5561
rect 296 5160 3464 5184
rect 296 2040 320 5160
rect 3440 2040 3464 5160
rect 296 2016 3464 2040
rect -498 1639 -178 1961
rect -4002 1560 -834 1584
rect -4002 -1560 -3978 1560
rect -858 -1560 -834 1560
rect -4002 -1584 -834 -1560
rect -4796 -1961 -4476 -1639
rect -8300 -2040 -5132 -2016
rect -8300 -5160 -8276 -2040
rect -5156 -5160 -5132 -2040
rect -8300 -5184 -5132 -5160
rect -6876 -5616 -6556 -5184
rect -4796 -5239 -4754 -1961
rect -4518 -5239 -4476 -1961
rect -2578 -2016 -2258 -1584
rect -498 -1639 -456 1639
rect -220 -1639 -178 1639
rect 1720 1584 2040 2016
rect 3800 1961 3842 5239
rect 4078 1961 4120 5239
rect 6018 5184 6338 5616
rect 8098 5561 8140 8839
rect 8376 5561 8418 8839
rect 8098 5239 8418 5561
rect 4594 5160 7762 5184
rect 4594 2040 4618 5160
rect 7738 2040 7762 5160
rect 4594 2016 7762 2040
rect 3800 1639 4120 1961
rect 296 1560 3464 1584
rect 296 -1560 320 1560
rect 3440 -1560 3464 1560
rect 296 -1584 3464 -1560
rect -498 -1961 -178 -1639
rect -4002 -2040 -834 -2016
rect -4002 -5160 -3978 -2040
rect -858 -5160 -834 -2040
rect -4002 -5184 -834 -5160
rect -4796 -5561 -4476 -5239
rect -8300 -5640 -5132 -5616
rect -8300 -8760 -8276 -5640
rect -5156 -8760 -5132 -5640
rect -8300 -8784 -5132 -8760
rect -6876 -9000 -6556 -8784
rect -4796 -8839 -4754 -5561
rect -4518 -8839 -4476 -5561
rect -2578 -5616 -2258 -5184
rect -498 -5239 -456 -1961
rect -220 -5239 -178 -1961
rect 1720 -2016 2040 -1584
rect 3800 -1639 3842 1639
rect 4078 -1639 4120 1639
rect 6018 1584 6338 2016
rect 8098 1961 8140 5239
rect 8376 1961 8418 5239
rect 8098 1639 8418 1961
rect 4594 1560 7762 1584
rect 4594 -1560 4618 1560
rect 7738 -1560 7762 1560
rect 4594 -1584 7762 -1560
rect 3800 -1961 4120 -1639
rect 296 -2040 3464 -2016
rect 296 -5160 320 -2040
rect 3440 -5160 3464 -2040
rect 296 -5184 3464 -5160
rect -498 -5561 -178 -5239
rect -4002 -5640 -834 -5616
rect -4002 -8760 -3978 -5640
rect -858 -8760 -834 -5640
rect -4002 -8784 -834 -8760
rect -4796 -9000 -4476 -8839
rect -2578 -9000 -2258 -8784
rect -498 -8839 -456 -5561
rect -220 -8839 -178 -5561
rect 1720 -5616 2040 -5184
rect 3800 -5239 3842 -1961
rect 4078 -5239 4120 -1961
rect 6018 -2016 6338 -1584
rect 8098 -1639 8140 1639
rect 8376 -1639 8418 1639
rect 8098 -1961 8418 -1639
rect 4594 -2040 7762 -2016
rect 4594 -5160 4618 -2040
rect 7738 -5160 7762 -2040
rect 4594 -5184 7762 -5160
rect 3800 -5561 4120 -5239
rect 296 -5640 3464 -5616
rect 296 -8760 320 -5640
rect 3440 -8760 3464 -5640
rect 296 -8784 3464 -8760
rect -498 -9000 -178 -8839
rect 1720 -9000 2040 -8784
rect 3800 -8839 3842 -5561
rect 4078 -8839 4120 -5561
rect 6018 -5616 6338 -5184
rect 8098 -5239 8140 -1961
rect 8376 -5239 8418 -1961
rect 8098 -5561 8418 -5239
rect 4594 -5640 7762 -5616
rect 4594 -8760 4618 -5640
rect 7738 -8760 7762 -5640
rect 4594 -8784 7762 -8760
rect 3800 -9000 4120 -8839
rect 6018 -9000 6338 -8784
rect 8098 -8839 8140 -5561
rect 8376 -8839 8418 -5561
rect 8098 -9000 8418 -8839
<< properties >>
string FIXED_BBOX 4498 5520 7858 8880
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 16.0 l 16.0 val 524.159 carea 2.00 cperi 0.19 nx 4 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
