magic
tech sky130A
magscale 1 2
timestamp 1717363523
<< nwell >>
rect -325 -1627 325 1627
<< pmos >>
rect -129 1208 -29 1408
rect 29 1208 129 1408
rect -129 772 -29 972
rect 29 772 129 972
rect -129 336 -29 536
rect 29 336 129 536
rect -129 -100 -29 100
rect 29 -100 129 100
rect -129 -536 -29 -336
rect 29 -536 129 -336
rect -129 -972 -29 -772
rect 29 -972 129 -772
rect -129 -1408 -29 -1208
rect 29 -1408 129 -1208
<< pdiff >>
rect -187 1396 -129 1408
rect -187 1220 -175 1396
rect -141 1220 -129 1396
rect -187 1208 -129 1220
rect -29 1396 29 1408
rect -29 1220 -17 1396
rect 17 1220 29 1396
rect -29 1208 29 1220
rect 129 1396 187 1408
rect 129 1220 141 1396
rect 175 1220 187 1396
rect 129 1208 187 1220
rect -187 960 -129 972
rect -187 784 -175 960
rect -141 784 -129 960
rect -187 772 -129 784
rect -29 960 29 972
rect -29 784 -17 960
rect 17 784 29 960
rect -29 772 29 784
rect 129 960 187 972
rect 129 784 141 960
rect 175 784 187 960
rect 129 772 187 784
rect -187 524 -129 536
rect -187 348 -175 524
rect -141 348 -129 524
rect -187 336 -129 348
rect -29 524 29 536
rect -29 348 -17 524
rect 17 348 29 524
rect -29 336 29 348
rect 129 524 187 536
rect 129 348 141 524
rect 175 348 187 524
rect 129 336 187 348
rect -187 88 -129 100
rect -187 -88 -175 88
rect -141 -88 -129 88
rect -187 -100 -129 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 129 88 187 100
rect 129 -88 141 88
rect 175 -88 187 88
rect 129 -100 187 -88
rect -187 -348 -129 -336
rect -187 -524 -175 -348
rect -141 -524 -129 -348
rect -187 -536 -129 -524
rect -29 -348 29 -336
rect -29 -524 -17 -348
rect 17 -524 29 -348
rect -29 -536 29 -524
rect 129 -348 187 -336
rect 129 -524 141 -348
rect 175 -524 187 -348
rect 129 -536 187 -524
rect -187 -784 -129 -772
rect -187 -960 -175 -784
rect -141 -960 -129 -784
rect -187 -972 -129 -960
rect -29 -784 29 -772
rect -29 -960 -17 -784
rect 17 -960 29 -784
rect -29 -972 29 -960
rect 129 -784 187 -772
rect 129 -960 141 -784
rect 175 -960 187 -784
rect 129 -972 187 -960
rect -187 -1220 -129 -1208
rect -187 -1396 -175 -1220
rect -141 -1396 -129 -1220
rect -187 -1408 -129 -1396
rect -29 -1220 29 -1208
rect -29 -1396 -17 -1220
rect 17 -1396 29 -1220
rect -29 -1408 29 -1396
rect 129 -1220 187 -1208
rect 129 -1396 141 -1220
rect 175 -1396 187 -1220
rect 129 -1408 187 -1396
<< pdiffc >>
rect -175 1220 -141 1396
rect -17 1220 17 1396
rect 141 1220 175 1396
rect -175 784 -141 960
rect -17 784 17 960
rect 141 784 175 960
rect -175 348 -141 524
rect -17 348 17 524
rect 141 348 175 524
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect -175 -524 -141 -348
rect -17 -524 17 -348
rect 141 -524 175 -348
rect -175 -960 -141 -784
rect -17 -960 17 -784
rect 141 -960 175 -784
rect -175 -1396 -141 -1220
rect -17 -1396 17 -1220
rect 141 -1396 175 -1220
<< nsubdiff >>
rect -289 1557 -193 1591
rect 193 1557 289 1591
rect -289 1495 -255 1557
rect 255 1495 289 1557
rect -289 -1557 -255 -1495
rect 255 -1557 289 -1495
rect -289 -1591 -193 -1557
rect 193 -1591 289 -1557
<< nsubdiffcont >>
rect -193 1557 193 1591
rect -289 -1495 -255 1495
rect 255 -1495 289 1495
rect -193 -1591 193 -1557
<< poly >>
rect -129 1489 -29 1505
rect -129 1455 -113 1489
rect -45 1455 -29 1489
rect -129 1408 -29 1455
rect 29 1489 129 1505
rect 29 1455 45 1489
rect 113 1455 129 1489
rect 29 1408 129 1455
rect -129 1161 -29 1208
rect -129 1127 -113 1161
rect -45 1127 -29 1161
rect -129 1111 -29 1127
rect 29 1161 129 1208
rect 29 1127 45 1161
rect 113 1127 129 1161
rect 29 1111 129 1127
rect -129 1053 -29 1069
rect -129 1019 -113 1053
rect -45 1019 -29 1053
rect -129 972 -29 1019
rect 29 1053 129 1069
rect 29 1019 45 1053
rect 113 1019 129 1053
rect 29 972 129 1019
rect -129 725 -29 772
rect -129 691 -113 725
rect -45 691 -29 725
rect -129 675 -29 691
rect 29 725 129 772
rect 29 691 45 725
rect 113 691 129 725
rect 29 675 129 691
rect -129 617 -29 633
rect -129 583 -113 617
rect -45 583 -29 617
rect -129 536 -29 583
rect 29 617 129 633
rect 29 583 45 617
rect 113 583 129 617
rect 29 536 129 583
rect -129 289 -29 336
rect -129 255 -113 289
rect -45 255 -29 289
rect -129 239 -29 255
rect 29 289 129 336
rect 29 255 45 289
rect 113 255 129 289
rect 29 239 129 255
rect -129 181 -29 197
rect -129 147 -113 181
rect -45 147 -29 181
rect -129 100 -29 147
rect 29 181 129 197
rect 29 147 45 181
rect 113 147 129 181
rect 29 100 129 147
rect -129 -147 -29 -100
rect -129 -181 -113 -147
rect -45 -181 -29 -147
rect -129 -197 -29 -181
rect 29 -147 129 -100
rect 29 -181 45 -147
rect 113 -181 129 -147
rect 29 -197 129 -181
rect -129 -255 -29 -239
rect -129 -289 -113 -255
rect -45 -289 -29 -255
rect -129 -336 -29 -289
rect 29 -255 129 -239
rect 29 -289 45 -255
rect 113 -289 129 -255
rect 29 -336 129 -289
rect -129 -583 -29 -536
rect -129 -617 -113 -583
rect -45 -617 -29 -583
rect -129 -633 -29 -617
rect 29 -583 129 -536
rect 29 -617 45 -583
rect 113 -617 129 -583
rect 29 -633 129 -617
rect -129 -691 -29 -675
rect -129 -725 -113 -691
rect -45 -725 -29 -691
rect -129 -772 -29 -725
rect 29 -691 129 -675
rect 29 -725 45 -691
rect 113 -725 129 -691
rect 29 -772 129 -725
rect -129 -1019 -29 -972
rect -129 -1053 -113 -1019
rect -45 -1053 -29 -1019
rect -129 -1069 -29 -1053
rect 29 -1019 129 -972
rect 29 -1053 45 -1019
rect 113 -1053 129 -1019
rect 29 -1069 129 -1053
rect -129 -1127 -29 -1111
rect -129 -1161 -113 -1127
rect -45 -1161 -29 -1127
rect -129 -1208 -29 -1161
rect 29 -1127 129 -1111
rect 29 -1161 45 -1127
rect 113 -1161 129 -1127
rect 29 -1208 129 -1161
rect -129 -1455 -29 -1408
rect -129 -1489 -113 -1455
rect -45 -1489 -29 -1455
rect -129 -1505 -29 -1489
rect 29 -1455 129 -1408
rect 29 -1489 45 -1455
rect 113 -1489 129 -1455
rect 29 -1505 129 -1489
<< polycont >>
rect -113 1455 -45 1489
rect 45 1455 113 1489
rect -113 1127 -45 1161
rect 45 1127 113 1161
rect -113 1019 -45 1053
rect 45 1019 113 1053
rect -113 691 -45 725
rect 45 691 113 725
rect -113 583 -45 617
rect 45 583 113 617
rect -113 255 -45 289
rect 45 255 113 289
rect -113 147 -45 181
rect 45 147 113 181
rect -113 -181 -45 -147
rect 45 -181 113 -147
rect -113 -289 -45 -255
rect 45 -289 113 -255
rect -113 -617 -45 -583
rect 45 -617 113 -583
rect -113 -725 -45 -691
rect 45 -725 113 -691
rect -113 -1053 -45 -1019
rect 45 -1053 113 -1019
rect -113 -1161 -45 -1127
rect 45 -1161 113 -1127
rect -113 -1489 -45 -1455
rect 45 -1489 113 -1455
<< locali >>
rect -289 1557 -193 1591
rect 193 1557 289 1591
rect -289 1495 -255 1557
rect 255 1495 289 1557
rect -129 1455 -113 1489
rect -45 1455 -29 1489
rect 29 1455 45 1489
rect 113 1455 129 1489
rect -175 1396 -141 1412
rect -175 1204 -141 1220
rect -17 1396 17 1412
rect -17 1204 17 1220
rect 141 1396 175 1412
rect 141 1204 175 1220
rect -129 1127 -113 1161
rect -45 1127 -29 1161
rect 29 1127 45 1161
rect 113 1127 129 1161
rect -129 1019 -113 1053
rect -45 1019 -29 1053
rect 29 1019 45 1053
rect 113 1019 129 1053
rect -175 960 -141 976
rect -175 768 -141 784
rect -17 960 17 976
rect -17 768 17 784
rect 141 960 175 976
rect 141 768 175 784
rect -129 691 -113 725
rect -45 691 -29 725
rect 29 691 45 725
rect 113 691 129 725
rect -129 583 -113 617
rect -45 583 -29 617
rect 29 583 45 617
rect 113 583 129 617
rect -175 524 -141 540
rect -175 332 -141 348
rect -17 524 17 540
rect -17 332 17 348
rect 141 524 175 540
rect 141 332 175 348
rect -129 255 -113 289
rect -45 255 -29 289
rect 29 255 45 289
rect 113 255 129 289
rect -129 147 -113 181
rect -45 147 -29 181
rect 29 147 45 181
rect 113 147 129 181
rect -175 88 -141 104
rect -175 -104 -141 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 141 88 175 104
rect 141 -104 175 -88
rect -129 -181 -113 -147
rect -45 -181 -29 -147
rect 29 -181 45 -147
rect 113 -181 129 -147
rect -129 -289 -113 -255
rect -45 -289 -29 -255
rect 29 -289 45 -255
rect 113 -289 129 -255
rect -175 -348 -141 -332
rect -175 -540 -141 -524
rect -17 -348 17 -332
rect -17 -540 17 -524
rect 141 -348 175 -332
rect 141 -540 175 -524
rect -129 -617 -113 -583
rect -45 -617 -29 -583
rect 29 -617 45 -583
rect 113 -617 129 -583
rect -129 -725 -113 -691
rect -45 -725 -29 -691
rect 29 -725 45 -691
rect 113 -725 129 -691
rect -175 -784 -141 -768
rect -175 -976 -141 -960
rect -17 -784 17 -768
rect -17 -976 17 -960
rect 141 -784 175 -768
rect 141 -976 175 -960
rect -129 -1053 -113 -1019
rect -45 -1053 -29 -1019
rect 29 -1053 45 -1019
rect 113 -1053 129 -1019
rect -129 -1161 -113 -1127
rect -45 -1161 -29 -1127
rect 29 -1161 45 -1127
rect 113 -1161 129 -1127
rect -175 -1220 -141 -1204
rect -175 -1412 -141 -1396
rect -17 -1220 17 -1204
rect -17 -1412 17 -1396
rect 141 -1220 175 -1204
rect 141 -1412 175 -1396
rect -129 -1489 -113 -1455
rect -45 -1489 -29 -1455
rect 29 -1489 45 -1455
rect 113 -1489 129 -1455
rect -289 -1557 -255 -1495
rect 255 -1557 289 -1495
rect -289 -1591 -193 -1557
rect 193 -1591 289 -1557
<< viali >>
rect -113 1455 -45 1489
rect 45 1455 113 1489
rect -175 1220 -141 1396
rect -17 1220 17 1396
rect 141 1220 175 1396
rect -113 1127 -45 1161
rect 45 1127 113 1161
rect -113 1019 -45 1053
rect 45 1019 113 1053
rect -175 784 -141 960
rect -17 784 17 960
rect 141 784 175 960
rect -113 691 -45 725
rect 45 691 113 725
rect -113 583 -45 617
rect 45 583 113 617
rect -175 348 -141 524
rect -17 348 17 524
rect 141 348 175 524
rect -113 255 -45 289
rect 45 255 113 289
rect -113 147 -45 181
rect 45 147 113 181
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect -113 -181 -45 -147
rect 45 -181 113 -147
rect -113 -289 -45 -255
rect 45 -289 113 -255
rect -175 -524 -141 -348
rect -17 -524 17 -348
rect 141 -524 175 -348
rect -113 -617 -45 -583
rect 45 -617 113 -583
rect -113 -725 -45 -691
rect 45 -725 113 -691
rect -175 -960 -141 -784
rect -17 -960 17 -784
rect 141 -960 175 -784
rect -113 -1053 -45 -1019
rect 45 -1053 113 -1019
rect -113 -1161 -45 -1127
rect 45 -1161 113 -1127
rect -175 -1396 -141 -1220
rect -17 -1396 17 -1220
rect 141 -1396 175 -1220
rect -113 -1489 -45 -1455
rect 45 -1489 113 -1455
<< metal1 >>
rect -125 1489 -33 1495
rect -125 1455 -113 1489
rect -45 1455 -33 1489
rect -125 1449 -33 1455
rect 33 1489 125 1495
rect 33 1455 45 1489
rect 113 1455 125 1489
rect 33 1449 125 1455
rect -181 1396 -135 1408
rect -181 1220 -175 1396
rect -141 1220 -135 1396
rect -181 1208 -135 1220
rect -23 1396 23 1408
rect -23 1220 -17 1396
rect 17 1220 23 1396
rect -23 1208 23 1220
rect 135 1396 181 1408
rect 135 1220 141 1396
rect 175 1220 181 1396
rect 135 1208 181 1220
rect -125 1161 -33 1167
rect -125 1127 -113 1161
rect -45 1127 -33 1161
rect -125 1121 -33 1127
rect 33 1161 125 1167
rect 33 1127 45 1161
rect 113 1127 125 1161
rect 33 1121 125 1127
rect -125 1053 -33 1059
rect -125 1019 -113 1053
rect -45 1019 -33 1053
rect -125 1013 -33 1019
rect 33 1053 125 1059
rect 33 1019 45 1053
rect 113 1019 125 1053
rect 33 1013 125 1019
rect -181 960 -135 972
rect -181 784 -175 960
rect -141 784 -135 960
rect -181 772 -135 784
rect -23 960 23 972
rect -23 784 -17 960
rect 17 784 23 960
rect -23 772 23 784
rect 135 960 181 972
rect 135 784 141 960
rect 175 784 181 960
rect 135 772 181 784
rect -125 725 -33 731
rect -125 691 -113 725
rect -45 691 -33 725
rect -125 685 -33 691
rect 33 725 125 731
rect 33 691 45 725
rect 113 691 125 725
rect 33 685 125 691
rect -125 617 -33 623
rect -125 583 -113 617
rect -45 583 -33 617
rect -125 577 -33 583
rect 33 617 125 623
rect 33 583 45 617
rect 113 583 125 617
rect 33 577 125 583
rect -181 524 -135 536
rect -181 348 -175 524
rect -141 348 -135 524
rect -181 336 -135 348
rect -23 524 23 536
rect -23 348 -17 524
rect 17 348 23 524
rect -23 336 23 348
rect 135 524 181 536
rect 135 348 141 524
rect 175 348 181 524
rect 135 336 181 348
rect -125 289 -33 295
rect -125 255 -113 289
rect -45 255 -33 289
rect -125 249 -33 255
rect 33 289 125 295
rect 33 255 45 289
rect 113 255 125 289
rect 33 249 125 255
rect -125 181 -33 187
rect -125 147 -113 181
rect -45 147 -33 181
rect -125 141 -33 147
rect 33 181 125 187
rect 33 147 45 181
rect 113 147 125 181
rect 33 141 125 147
rect -181 88 -135 100
rect -181 -88 -175 88
rect -141 -88 -135 88
rect -181 -100 -135 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 135 88 181 100
rect 135 -88 141 88
rect 175 -88 181 88
rect 135 -100 181 -88
rect -125 -147 -33 -141
rect -125 -181 -113 -147
rect -45 -181 -33 -147
rect -125 -187 -33 -181
rect 33 -147 125 -141
rect 33 -181 45 -147
rect 113 -181 125 -147
rect 33 -187 125 -181
rect -125 -255 -33 -249
rect -125 -289 -113 -255
rect -45 -289 -33 -255
rect -125 -295 -33 -289
rect 33 -255 125 -249
rect 33 -289 45 -255
rect 113 -289 125 -255
rect 33 -295 125 -289
rect -181 -348 -135 -336
rect -181 -524 -175 -348
rect -141 -524 -135 -348
rect -181 -536 -135 -524
rect -23 -348 23 -336
rect -23 -524 -17 -348
rect 17 -524 23 -348
rect -23 -536 23 -524
rect 135 -348 181 -336
rect 135 -524 141 -348
rect 175 -524 181 -348
rect 135 -536 181 -524
rect -125 -583 -33 -577
rect -125 -617 -113 -583
rect -45 -617 -33 -583
rect -125 -623 -33 -617
rect 33 -583 125 -577
rect 33 -617 45 -583
rect 113 -617 125 -583
rect 33 -623 125 -617
rect -125 -691 -33 -685
rect -125 -725 -113 -691
rect -45 -725 -33 -691
rect -125 -731 -33 -725
rect 33 -691 125 -685
rect 33 -725 45 -691
rect 113 -725 125 -691
rect 33 -731 125 -725
rect -181 -784 -135 -772
rect -181 -960 -175 -784
rect -141 -960 -135 -784
rect -181 -972 -135 -960
rect -23 -784 23 -772
rect -23 -960 -17 -784
rect 17 -960 23 -784
rect -23 -972 23 -960
rect 135 -784 181 -772
rect 135 -960 141 -784
rect 175 -960 181 -784
rect 135 -972 181 -960
rect -125 -1019 -33 -1013
rect -125 -1053 -113 -1019
rect -45 -1053 -33 -1019
rect -125 -1059 -33 -1053
rect 33 -1019 125 -1013
rect 33 -1053 45 -1019
rect 113 -1053 125 -1019
rect 33 -1059 125 -1053
rect -125 -1127 -33 -1121
rect -125 -1161 -113 -1127
rect -45 -1161 -33 -1127
rect -125 -1167 -33 -1161
rect 33 -1127 125 -1121
rect 33 -1161 45 -1127
rect 113 -1161 125 -1127
rect 33 -1167 125 -1161
rect -181 -1220 -135 -1208
rect -181 -1396 -175 -1220
rect -141 -1396 -135 -1220
rect -181 -1408 -135 -1396
rect -23 -1220 23 -1208
rect -23 -1396 -17 -1220
rect 17 -1396 23 -1220
rect -23 -1408 23 -1396
rect 135 -1220 181 -1208
rect 135 -1396 141 -1220
rect 175 -1396 181 -1220
rect 135 -1408 181 -1396
rect -125 -1455 -33 -1449
rect -125 -1489 -113 -1455
rect -45 -1489 -33 -1455
rect -125 -1495 -33 -1489
rect 33 -1455 125 -1449
rect 33 -1489 45 -1455
rect 113 -1489 125 -1455
rect 33 -1495 125 -1489
<< properties >>
string FIXED_BBOX -272 -1574 272 1574
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 0.5 m 7 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
