** sch_path: /home/cmos/Downloads/sky130_ef_ip__bgrref_por/cace/startup_sim.sch
**.subckt startup_sim por porb porb_h
*.opin por
*.opin porb
*.opin porb_h
XDUT vbg por avss avdd dvdd porb dvss porb_h VCC VSS sky130_ef_ip__bgrref_por W_N=1 L_N=0.2 W_P=1
+ L_P=0.2 m=1
Vdvss dvss GND DC {Vdvss}
Vavdd avdd GND PULSE 0 {Vavdd} 10e-9 1e-3 1e-3 100e-3 200e-3
Vavss avss GND DC {Vavss}
Vdvdd dvdd GND PULSE 0 {Vdvdd} 10e-9 1.1e-3 1e-3 200e-3 400e-3
Vvbg vbg GND PULSE 0 {Vvbg} 10e-9 0.5e-3 1e-3 200e-3 400e-3
**** begin user architecture code


* CACE gensim simulation file {filename}
* Generated by CACE gensim, Efabless Corporation (c) 2024
* Find the powerup simulation of POR

.include {DUT_path}
.include {PDK_ROOT}/{PDK}/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice
.include {PDK_ROOT}/{PDK}/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

.lib {PDK_ROOT}/{PDK}/libs.tech/combined/sky130.lib.spice {corner}

.option TEMP={temperature}
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1




.control
save all
tran .1u 2m
*plot AVDD por porb+6.8 porb_h+3.4
wrdata {simpath}/{filename}_{N}.data V(por) V(porb) V(porb_h) V(avdd) V(bg) V(dvdd)

quit
.endc


**** end user architecture code
**.ends

* expanding   symbol:  sky130_ef_ip__bgrref_por.sym # of pins=8
** sym_path: /home/cmos/Downloads/sky130_ef_ip__bgrref_por/xschem/sky130_ef_ip__bgrref_por.sym
** sch_path: /home/cmos/Downloads/sky130_ef_ip__bgrref_por/xschem/sky130_ef_ip__bgrref_por.sch
.subckt sky130_ef_ip__bgrref_por vbg por avss avdd dvdd porb dvss porb_h VCCBPIN VSSBPIN  W_N=1 L_N=0.2 W_P=1 L_P=0.2
*.iopin avdd
*.opin por
*.iopin avss
*.iopin dvdd
*.opin porb
*.ipin vbg
*.opin porb_h
*.iopin dvss
XM1 avdd avdd net3 avss sky130_fd_pr__nfet_05v0_nvt L=0.9 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf
+ * 0.29' as='int((nf+2)/2) * W / nf * 0.29' pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2)
+ * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2 m=2
Vr1 net3 net1 0
.save i(vr1)
E1 vindiff GND Vinp Vinn 1
x1 Iref Vinn Vinp RST avss avdd dvdd comparator
XR1 avss Vinn avss sky130_fd_pr__res_xhigh_po_0p35 L=235 mult=1 m=1
XR10 Vinn Vinp avss sky130_fd_pr__res_xhigh_po_0p35 L=10.4 mult=1 m=1
XR12 Vinp net1 avss sky130_fd_pr__res_xhigh_po_0p35 L=120 mult=1 m=1
x2 RST por dvdd dvss vbg avdd porb porb_h net2 delayPulse
Vr2 net2 Iref 0
.save i(vr2)
.ends


* expanding   symbol:  comparator.sym # of pins=7
** sym_path: /home/cmos/Downloads/sky130_ef_ip__bgrref_por/xschem/comparator.sym
** sch_path: /home/cmos/Downloads/sky130_ef_ip__bgrref_por/xschem/comparator.sch
.subckt comparator Iref Vinn Vinp RST VSS AVDD DVDD
*.ipin AVDD
*.opin RST
*.ipin VSS
*.iopin Iref
*.ipin Vinn
*.ipin Vinp
*.ipin DVDD
v1 AVDD net3 0
.save i(v1)
v2 AVDD net4 0
.save i(v2)
XM1 net5 vbn VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM3 vbp vbp net3 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=24 m=24
XM2 vt vbp net4 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=24 m=24
v4 net6 vo1 0
.save i(v4)
XM9 VD Vinn VS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM10 net1 Vinp VS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM5 Iref Iref VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM7 vo vt AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
v3 VS net5 0
.save i(v3)
XM11 VD Vinn VY VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6
x1 VD VS VY AVDD VSS Sel mux2to1
XM6 vo vbn VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6
v6 net7 net2 0
.save i(v6)
XM14 vo1 vo VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15 net6 vo DVDD DVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 net2 vo1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13 net7 vo1 DVDD DVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x2 vo1 Sel DVDD VSS AVDD levelShifter
v5 net8 RST 0
.save i(v5)
XM16 RST net2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM17 net8 net2 DVDD DVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XC1 vbn VSS sky130_fd_pr__cap_mim_m3_2 W=11 L=11 MF=1 m=1
XM4 vbp vbp net1 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=16 m=16
XM8 vt vt VD VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=16 m=16
XR9 Iref vbn VSS sky130_fd_pr__res_xhigh_po W=1 L=300 mult=1 m=1
.ends


* expanding   symbol:  delayPulse.sym # of pins=9
** sym_path: /home/cmos/Downloads/sky130_ef_ip__bgrref_por/xschem/delayPulse.sym
** sch_path: /home/cmos/Downloads/sky130_ef_ip__bgrref_por/xschem/delayPulse.sch
.subckt delayPulse din por VCCL VSS Vbg VCCH porb porb_h Iref
*.ipin VCCL
*.ipin VSS
*.ipin din
*.ipin Vbg
*.opin por
*.ipin VCCH
*.opin porb
*.opin porb_h
*.iopin Iref
v9 net20 VT2 0
.save i(v9)
v1 net21 Td_S 0
.save i(v1)
v3 net22 net1 0
.save i(v3)
x1 Td_L Td_Sd VSS VSS VCCL VCCL outxor sky130_fd_sc_hd__xor2_1
x3 porb porb_h VCCL VSS VCCH levelShifter
XM2 net22 din VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM3 net21 net1 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM5 VT2 net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 net1 din VSS VSS sky130_fd_pr__nfet_01v8 L=0.3 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM8 Td_S net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.3 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM10 net20 net1 net13 VCCL sky130_fd_pr__pfet_01v8 L=0.3 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
v5 net23 VT3 0
.save i(v5)
v6 net24 net4 0
.save i(v6)
XM13 net4 VT3 VSS VSS sky130_fd_pr__nfet_01v8 L=0.3 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM14 net24 VT3 net5 net5 sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
x4 net2 VSS VCCL TieH_1p8
v2 net11 Iref 0
.save i(v2)
XM11 vbn1 net8 net6 VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM17 vbp2 vbn1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM18 net6 net7 VCCH VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM19 vbn1 vbn1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=14 nf=7 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM24 net8 net8 net7 VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM25 net7 net7 VCCH VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=16 nf=8 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM26 net19 Vbg net9 VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM28 net10 net7 VCCH VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM6 VT3 VT2 net3 VSS sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 net23 VT2 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.3 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 vbp2 vbp2 vbp1 VCCL sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15 vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=7 m=7
XM16 net12 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM20 net13 vbp2 net12 VCCL sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM21 net3 vbn1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM22 net14 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM23 net5 vbp2 net14 VCCL sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM27 net15 net4 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM29 net15 net4 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM30 Td_L net15 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM31 Td_L net15 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM32 net16 Td_S VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM33 net16 Td_S VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM34 net17 net16 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM35 net17 net16 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM36 Td_Sd net18 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM38 net18 net17 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM39 net18 net17 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x6 outxor VSS VSS VCCL VCCL rstn sky130_fd_sc_hvl__buf_8
XC4 net17 VSS sky130_fd_pr__cap_mim_m3_2 W=10 L=10 MF=2 m=2
XC7 VT2 VSS sky130_fd_pr__cap_mim_m3_2 W=16 L=16 MF=40 m=40
XC2 VT3 VSS sky130_fd_pr__cap_mim_m3_2 W=16 L=16 MF=40 m=40
XC8 net16 VSS sky130_fd_pr__cap_mim_m3_2 W=10 L=10 MF=2 m=2
XC9 net18 VSS sky130_fd_pr__cap_mim_m3_2 W=10 L=10 MF=2 m=2
XM40 Td_Sd net18 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM37 net11 net8 net10 VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
v4 net8 net19 0
.save i(v4)
x5 rstn net2 Td_S VSS VSS VCCL VCCL porb sky130_fd_sc_hd__dfrtn_1
x2 Td_S net2 Td_Lb VSS VSS VCCL VCCL por sky130_fd_sc_hd__dfrtp_1
XM4 Td_Lb Td_L VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM9 Td_Lb Td_L VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XC1 vbn1 VSS sky130_fd_pr__cap_mim_m3_2 W=16 L=16 MF=2 m=2
XC5 VCCH net7 sky130_fd_pr__cap_mim_m3_2 W=16 L=16 MF=2 m=2
XC6 VCCL vbp1 sky130_fd_pr__cap_mim_m3_2 W=16 L=16 MF=2 m=2
XC3 VCCH net8 sky130_fd_pr__cap_mim_m3_2 W=8 L=8 MF=2 m=2
XR9 net25 net9 VSS sky130_fd_pr__res_xhigh_po W=1 L=350 mult=1 m=1
XR6 VSS net25 VSS sky130_fd_pr__res_xhigh_po W=1 L=350 mult=1 m=1
.ends


* expanding   symbol:  mux2to1.sym # of pins=6
** sym_path: /home/cmos/Downloads/sky130_ef_ip__bgrref_por/xschem/mux2to1.sym
** sch_path: /home/cmos/Downloads/sky130_ef_ip__bgrref_por/xschem/mux2to1.sch
.subckt mux2to1 A1 A0 Z VCC VSS S
*.ipin VCC
*.ipin VSS
*.ipin A0
*.ipin A1
*.iopin Z
*.ipin S
x2 Z A0 S SB VCC VSS passgate_3p3 W_N=1 L_N=0.2 W_P=1 L_P=0.2 m=1
x1 Z A1 SB S VCC VSS passgate_3p3 W_N=1 L_N=0.2 W_P=1 L_P=0.2 m=1
XM12 SB S VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
v9 net1 SB 0
.save i(v9)
XM13 net1 S VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  levelShifter.sym # of pins=5
** sym_path: /home/cmos/Downloads/sky130_ef_ip__bgrref_por/xschem/levelShifter.sym
** sch_path: /home/cmos/Downloads/sky130_ef_ip__bgrref_por/xschem/levelShifter.sch
.subckt levelShifter ain aout VCCL VSS VCCH
*.ipin VCCL
*.ipin VSS
*.ipin ain
*.opin aout
*.ipin VCCH
v6 net3 net2 0
.save i(v6)
XM12 net1 S1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM13 net3 net1 VCCH VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2.9 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
v5 net4 S1 0
.save i(v5)
XM6 S1 ain VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 net4 ain VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
v1 net5 net1 0
.save i(v1)
XM2 net5 net2 VCCH VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2.9 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM3 net2 S1B VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
v2 net6 S1B 0
.save i(v2)
XM4 S1B S1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net6 S1 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 aout net2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM8 aout net2 VCCH VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2.9 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
.ends


* expanding   symbol:  TieH_1p8.sym # of pins=3
** sym_path: /home/cmos/Downloads/sky130_ef_ip__bgrref_por/xschem/TieH_1p8.sym
** sch_path: /home/cmos/Downloads/sky130_ef_ip__bgrref_por/xschem/TieH_1p8.sch
.subckt TieH_1p8 TieH VSS VCC
*.ipin VCC
*.ipin VSS
*.iopin TieH
v2 net2 TieH 0
.save i(v2)
XM4 net1 net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net2 net1 VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  passgate_3p3.sym # of pins=4
** sym_path: /home/cmos/Downloads/sky130_ef_ip__bgrref_por/xschem/passgate_3p3.sym
** sch_path: /home/cmos/Downloads/sky130_ef_ip__bgrref_por/xschem/passgate_3p3.sch
.subckt passgate_3p3 Z A GP GN VCCBPIN VSSBPIN  W_N=1 L_N=0.2 W_P=1 L_P=0.2
*.iopin A
*.iopin Z
*.ipin GP
*.ipin GN
* noconn VCCBPIN
* noconn VSSBPIN
XM3 Z GP A VCCBPIN sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM4 Z GN A VSSBPIN sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 /
+ W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
