magic
tech sky130A
magscale 1 2
timestamp 1717363523
<< pwell >>
rect -201 -3382 201 3382
<< psubdiff >>
rect -165 3312 -69 3346
rect 69 3312 165 3346
rect -165 3250 -131 3312
rect 131 3250 165 3312
rect -165 -3312 -131 -3250
rect 131 -3312 165 -3250
rect -165 -3346 -69 -3312
rect 69 -3346 165 -3312
<< psubdiffcont >>
rect -69 3312 69 3346
rect -165 -3250 -131 3250
rect 131 -3250 165 3250
rect -69 -3346 69 -3312
<< xpolycontact >>
rect -35 2784 35 3216
rect -35 -3216 35 -2784
<< xpolyres >>
rect -35 -2784 35 2784
<< locali >>
rect -165 3312 -69 3346
rect 69 3312 165 3346
rect -165 3250 -131 3312
rect 131 3250 165 3312
rect -165 -3312 -131 -3250
rect 131 -3312 165 -3250
rect -165 -3346 -69 -3312
rect 69 -3346 165 -3312
<< viali >>
rect -19 2801 19 3198
rect -19 -3198 19 -2801
<< metal1 >>
rect -25 3198 25 3210
rect -25 2801 -19 3198
rect 19 2801 25 3198
rect -25 2789 25 2801
rect -25 -2801 25 -2789
rect -25 -3198 -19 -2801
rect 19 -3198 25 -2801
rect -25 -3210 25 -3198
<< properties >>
string FIXED_BBOX -148 -3329 148 3329
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 28.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 161.075k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
