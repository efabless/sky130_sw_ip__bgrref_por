magic
tech sky130A
magscale 1 2
timestamp 1718283729
<< pwell >>
rect -2926 -1582 2926 1582
<< psubdiff >>
rect -2890 1512 -2794 1546
rect 2794 1512 2890 1546
rect -2890 1450 -2856 1512
rect 2856 1450 2890 1512
rect -2890 -1512 -2856 -1450
rect 2856 -1512 2890 -1450
rect -2890 -1546 -2794 -1512
rect 2794 -1546 2890 -1512
<< psubdiffcont >>
rect -2794 1512 2794 1546
rect -2890 -1450 -2856 1450
rect 2856 -1450 2890 1450
rect -2794 -1546 2794 -1512
<< xpolycontact >>
rect -2760 984 -2622 1416
rect -2760 -1416 -2622 -984
rect -2526 984 -2388 1416
rect -2526 -1416 -2388 -984
rect -2292 984 -2154 1416
rect -2292 -1416 -2154 -984
rect -2058 984 -1920 1416
rect -2058 -1416 -1920 -984
rect -1824 984 -1686 1416
rect -1824 -1416 -1686 -984
rect -1590 984 -1452 1416
rect -1590 -1416 -1452 -984
rect -1356 984 -1218 1416
rect -1356 -1416 -1218 -984
rect -1122 984 -984 1416
rect -1122 -1416 -984 -984
rect -888 984 -750 1416
rect -888 -1416 -750 -984
rect -654 984 -516 1416
rect -654 -1416 -516 -984
rect -420 984 -282 1416
rect -420 -1416 -282 -984
rect -186 984 -48 1416
rect -186 -1416 -48 -984
rect 48 984 186 1416
rect 48 -1416 186 -984
rect 282 984 420 1416
rect 282 -1416 420 -984
rect 516 984 654 1416
rect 516 -1416 654 -984
rect 750 984 888 1416
rect 750 -1416 888 -984
rect 984 984 1122 1416
rect 984 -1416 1122 -984
rect 1218 984 1356 1416
rect 1218 -1416 1356 -984
rect 1452 984 1590 1416
rect 1452 -1416 1590 -984
rect 1686 984 1824 1416
rect 1686 -1416 1824 -984
rect 1920 984 2058 1416
rect 1920 -1416 2058 -984
rect 2154 984 2292 1416
rect 2154 -1416 2292 -984
rect 2388 984 2526 1416
rect 2388 -1416 2526 -984
rect 2622 984 2760 1416
rect 2622 -1416 2760 -984
<< xpolyres >>
rect -2760 -984 -2622 984
rect -2526 -984 -2388 984
rect -2292 -984 -2154 984
rect -2058 -984 -1920 984
rect -1824 -984 -1686 984
rect -1590 -984 -1452 984
rect -1356 -984 -1218 984
rect -1122 -984 -984 984
rect -888 -984 -750 984
rect -654 -984 -516 984
rect -420 -984 -282 984
rect -186 -984 -48 984
rect 48 -984 186 984
rect 282 -984 420 984
rect 516 -984 654 984
rect 750 -984 888 984
rect 984 -984 1122 984
rect 1218 -984 1356 984
rect 1452 -984 1590 984
rect 1686 -984 1824 984
rect 1920 -984 2058 984
rect 2154 -984 2292 984
rect 2388 -984 2526 984
rect 2622 -984 2760 984
<< locali >>
rect -2890 1512 -2794 1546
rect 2794 1512 2890 1546
rect -2890 1450 -2856 1512
rect 2856 1450 2890 1512
rect -2890 -1512 -2856 -1450
rect 2856 -1512 2890 -1450
rect -2890 -1546 -2794 -1512
rect 2794 -1546 2890 -1512
<< viali >>
rect -2744 1001 -2638 1398
rect -2510 1001 -2404 1398
rect -2276 1001 -2170 1398
rect -2042 1001 -1936 1398
rect -1808 1001 -1702 1398
rect -1574 1001 -1468 1398
rect -1340 1001 -1234 1398
rect -1106 1001 -1000 1398
rect -872 1001 -766 1398
rect -638 1001 -532 1398
rect -404 1001 -298 1398
rect -170 1001 -64 1398
rect 64 1001 170 1398
rect 298 1001 404 1398
rect 532 1001 638 1398
rect 766 1001 872 1398
rect 1000 1001 1106 1398
rect 1234 1001 1340 1398
rect 1468 1001 1574 1398
rect 1702 1001 1808 1398
rect 1936 1001 2042 1398
rect 2170 1001 2276 1398
rect 2404 1001 2510 1398
rect 2638 1001 2744 1398
rect -2744 -1398 -2638 -1001
rect -2510 -1398 -2404 -1001
rect -2276 -1398 -2170 -1001
rect -2042 -1398 -1936 -1001
rect -1808 -1398 -1702 -1001
rect -1574 -1398 -1468 -1001
rect -1340 -1398 -1234 -1001
rect -1106 -1398 -1000 -1001
rect -872 -1398 -766 -1001
rect -638 -1398 -532 -1001
rect -404 -1398 -298 -1001
rect -170 -1398 -64 -1001
rect 64 -1398 170 -1001
rect 298 -1398 404 -1001
rect 532 -1398 638 -1001
rect 766 -1398 872 -1001
rect 1000 -1398 1106 -1001
rect 1234 -1398 1340 -1001
rect 1468 -1398 1574 -1001
rect 1702 -1398 1808 -1001
rect 1936 -1398 2042 -1001
rect 2170 -1398 2276 -1001
rect 2404 -1398 2510 -1001
rect 2638 -1398 2744 -1001
<< metal1 >>
rect -2750 1398 -2632 1410
rect -2750 1001 -2744 1398
rect -2638 1001 -2632 1398
rect -2750 989 -2632 1001
rect -2516 1398 -2398 1410
rect -2516 1001 -2510 1398
rect -2404 1001 -2398 1398
rect -2516 989 -2398 1001
rect -2282 1398 -2164 1410
rect -2282 1001 -2276 1398
rect -2170 1001 -2164 1398
rect -2282 989 -2164 1001
rect -2048 1398 -1930 1410
rect -2048 1001 -2042 1398
rect -1936 1001 -1930 1398
rect -2048 989 -1930 1001
rect -1814 1398 -1696 1410
rect -1814 1001 -1808 1398
rect -1702 1001 -1696 1398
rect -1814 989 -1696 1001
rect -1580 1398 -1462 1410
rect -1580 1001 -1574 1398
rect -1468 1001 -1462 1398
rect -1580 989 -1462 1001
rect -1346 1398 -1228 1410
rect -1346 1001 -1340 1398
rect -1234 1001 -1228 1398
rect -1346 989 -1228 1001
rect -1112 1398 -994 1410
rect -1112 1001 -1106 1398
rect -1000 1001 -994 1398
rect -1112 989 -994 1001
rect -878 1398 -760 1410
rect -878 1001 -872 1398
rect -766 1001 -760 1398
rect -878 989 -760 1001
rect -644 1398 -526 1410
rect -644 1001 -638 1398
rect -532 1001 -526 1398
rect -644 989 -526 1001
rect -410 1398 -292 1410
rect -410 1001 -404 1398
rect -298 1001 -292 1398
rect -410 989 -292 1001
rect -176 1398 -58 1410
rect -176 1001 -170 1398
rect -64 1001 -58 1398
rect -176 989 -58 1001
rect 58 1398 176 1410
rect 58 1001 64 1398
rect 170 1001 176 1398
rect 58 989 176 1001
rect 292 1398 410 1410
rect 292 1001 298 1398
rect 404 1001 410 1398
rect 292 989 410 1001
rect 526 1398 644 1410
rect 526 1001 532 1398
rect 638 1001 644 1398
rect 526 989 644 1001
rect 760 1398 878 1410
rect 760 1001 766 1398
rect 872 1001 878 1398
rect 760 989 878 1001
rect 994 1398 1112 1410
rect 994 1001 1000 1398
rect 1106 1001 1112 1398
rect 994 989 1112 1001
rect 1228 1398 1346 1410
rect 1228 1001 1234 1398
rect 1340 1001 1346 1398
rect 1228 989 1346 1001
rect 1462 1398 1580 1410
rect 1462 1001 1468 1398
rect 1574 1001 1580 1398
rect 1462 989 1580 1001
rect 1696 1398 1814 1410
rect 1696 1001 1702 1398
rect 1808 1001 1814 1398
rect 1696 989 1814 1001
rect 1930 1398 2048 1410
rect 1930 1001 1936 1398
rect 2042 1001 2048 1398
rect 1930 989 2048 1001
rect 2164 1398 2282 1410
rect 2164 1001 2170 1398
rect 2276 1001 2282 1398
rect 2164 989 2282 1001
rect 2398 1398 2516 1410
rect 2398 1001 2404 1398
rect 2510 1001 2516 1398
rect 2398 989 2516 1001
rect 2632 1398 2750 1410
rect 2632 1001 2638 1398
rect 2744 1001 2750 1398
rect 2632 989 2750 1001
rect -2750 -1001 -2632 -989
rect -2750 -1398 -2744 -1001
rect -2638 -1398 -2632 -1001
rect -2750 -1410 -2632 -1398
rect -2516 -1001 -2398 -989
rect -2516 -1398 -2510 -1001
rect -2404 -1398 -2398 -1001
rect -2516 -1410 -2398 -1398
rect -2282 -1001 -2164 -989
rect -2282 -1398 -2276 -1001
rect -2170 -1398 -2164 -1001
rect -2282 -1410 -2164 -1398
rect -2048 -1001 -1930 -989
rect -2048 -1398 -2042 -1001
rect -1936 -1398 -1930 -1001
rect -2048 -1410 -1930 -1398
rect -1814 -1001 -1696 -989
rect -1814 -1398 -1808 -1001
rect -1702 -1398 -1696 -1001
rect -1814 -1410 -1696 -1398
rect -1580 -1001 -1462 -989
rect -1580 -1398 -1574 -1001
rect -1468 -1398 -1462 -1001
rect -1580 -1410 -1462 -1398
rect -1346 -1001 -1228 -989
rect -1346 -1398 -1340 -1001
rect -1234 -1398 -1228 -1001
rect -1346 -1410 -1228 -1398
rect -1112 -1001 -994 -989
rect -1112 -1398 -1106 -1001
rect -1000 -1398 -994 -1001
rect -1112 -1410 -994 -1398
rect -878 -1001 -760 -989
rect -878 -1398 -872 -1001
rect -766 -1398 -760 -1001
rect -878 -1410 -760 -1398
rect -644 -1001 -526 -989
rect -644 -1398 -638 -1001
rect -532 -1398 -526 -1001
rect -644 -1410 -526 -1398
rect -410 -1001 -292 -989
rect -410 -1398 -404 -1001
rect -298 -1398 -292 -1001
rect -410 -1410 -292 -1398
rect -176 -1001 -58 -989
rect -176 -1398 -170 -1001
rect -64 -1398 -58 -1001
rect -176 -1410 -58 -1398
rect 58 -1001 176 -989
rect 58 -1398 64 -1001
rect 170 -1398 176 -1001
rect 58 -1410 176 -1398
rect 292 -1001 410 -989
rect 292 -1398 298 -1001
rect 404 -1398 410 -1001
rect 292 -1410 410 -1398
rect 526 -1001 644 -989
rect 526 -1398 532 -1001
rect 638 -1398 644 -1001
rect 526 -1410 644 -1398
rect 760 -1001 878 -989
rect 760 -1398 766 -1001
rect 872 -1398 878 -1001
rect 760 -1410 878 -1398
rect 994 -1001 1112 -989
rect 994 -1398 1000 -1001
rect 1106 -1398 1112 -1001
rect 994 -1410 1112 -1398
rect 1228 -1001 1346 -989
rect 1228 -1398 1234 -1001
rect 1340 -1398 1346 -1001
rect 1228 -1410 1346 -1398
rect 1462 -1001 1580 -989
rect 1462 -1398 1468 -1001
rect 1574 -1398 1580 -1001
rect 1462 -1410 1580 -1398
rect 1696 -1001 1814 -989
rect 1696 -1398 1702 -1001
rect 1808 -1398 1814 -1001
rect 1696 -1410 1814 -1398
rect 1930 -1001 2048 -989
rect 1930 -1398 1936 -1001
rect 2042 -1398 2048 -1001
rect 1930 -1410 2048 -1398
rect 2164 -1001 2282 -989
rect 2164 -1398 2170 -1001
rect 2276 -1398 2282 -1001
rect 2164 -1410 2282 -1398
rect 2398 -1001 2516 -989
rect 2398 -1398 2404 -1001
rect 2510 -1398 2516 -1001
rect 2398 -1410 2516 -1398
rect 2632 -1001 2750 -989
rect 2632 -1398 2638 -1001
rect 2744 -1398 2750 -1001
rect 2632 -1410 2750 -1398
<< properties >>
string FIXED_BBOX -2873 -1529 2873 1529
string gencell sky130_fd_pr__res_xhigh_po_0p69
string library sky130
string parameters w 0.690 l 10 m 1 nx 24 wmin 0.690 lmin 0.50 rho 2000 val 29.531k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.690 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
