magic
tech sky130A
magscale 1 2
timestamp 1731450921
<< pwell >>
rect -450 -4182 450 4182
<< psubdiff >>
rect -414 4112 -318 4146
rect 318 4112 414 4146
rect -414 4050 -380 4112
rect 380 4050 414 4112
rect -414 -4112 -380 -4050
rect 380 -4112 414 -4050
rect -414 -4146 -318 -4112
rect 318 -4146 414 -4112
<< psubdiffcont >>
rect -318 4112 318 4146
rect -414 -4050 -380 4050
rect 380 -4050 414 4050
rect -318 -4146 318 -4112
<< xpolycontact >>
rect -284 3584 -214 4016
rect -284 -4016 -214 -3584
rect -118 3584 -48 4016
rect -118 -4016 -48 -3584
rect 48 3584 118 4016
rect 48 -4016 118 -3584
rect 214 3584 284 4016
rect 214 -4016 284 -3584
<< xpolyres >>
rect -284 -3584 -214 3584
rect -118 -3584 -48 3584
rect 48 -3584 118 3584
rect 214 -3584 284 3584
<< locali >>
rect -414 4112 -318 4146
rect 318 4112 414 4146
rect -414 4050 -380 4112
rect 380 4050 414 4112
rect -414 -4112 -380 -4050
rect 380 -4112 414 -4050
rect -414 -4146 -318 -4112
rect 318 -4146 414 -4112
<< viali >>
rect -268 3601 -230 3998
rect -102 3601 -64 3998
rect 64 3601 102 3998
rect 230 3601 268 3998
rect -268 -3998 -230 -3601
rect -102 -3998 -64 -3601
rect 64 -3998 102 -3601
rect 230 -3998 268 -3601
<< metal1 >>
rect -274 3998 -224 4010
rect -274 3601 -268 3998
rect -230 3601 -224 3998
rect -274 3589 -224 3601
rect -108 3998 -58 4010
rect -108 3601 -102 3998
rect -64 3601 -58 3998
rect -108 3589 -58 3601
rect 58 3998 108 4010
rect 58 3601 64 3998
rect 102 3601 108 3998
rect 58 3589 108 3601
rect 224 3998 274 4010
rect 224 3601 230 3998
rect 268 3601 274 3998
rect 224 3589 274 3601
rect -274 -3601 -224 -3589
rect -274 -3998 -268 -3601
rect -230 -3998 -224 -3601
rect -274 -4010 -224 -3998
rect -108 -3601 -58 -3589
rect -108 -3998 -102 -3601
rect -64 -3998 -58 -3601
rect -108 -4010 -58 -3998
rect 58 -3601 108 -3589
rect 58 -3998 64 -3601
rect 102 -3998 108 -3601
rect 58 -4010 108 -3998
rect 224 -3601 274 -3589
rect 224 -3998 230 -3601
rect 268 -3998 274 -3601
rect 224 -4010 274 -3998
<< properties >>
string FIXED_BBOX -397 -4129 397 4129
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 36 m 1 nx 4 wmin 0.350 lmin 0.50 class resistor rho 2000 val 206.789k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
