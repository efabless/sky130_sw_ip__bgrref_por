magic
tech sky130A
magscale 1 2
timestamp 1717363523
<< pwell >>
rect -308 -1385 308 1385
<< mvnmos >>
rect -80 727 80 1127
rect -80 109 80 509
rect -80 -509 80 -109
rect -80 -1127 80 -727
<< mvndiff >>
rect -138 1115 -80 1127
rect -138 739 -126 1115
rect -92 739 -80 1115
rect -138 727 -80 739
rect 80 1115 138 1127
rect 80 739 92 1115
rect 126 739 138 1115
rect 80 727 138 739
rect -138 497 -80 509
rect -138 121 -126 497
rect -92 121 -80 497
rect -138 109 -80 121
rect 80 497 138 509
rect 80 121 92 497
rect 126 121 138 497
rect 80 109 138 121
rect -138 -121 -80 -109
rect -138 -497 -126 -121
rect -92 -497 -80 -121
rect -138 -509 -80 -497
rect 80 -121 138 -109
rect 80 -497 92 -121
rect 126 -497 138 -121
rect 80 -509 138 -497
rect -138 -739 -80 -727
rect -138 -1115 -126 -739
rect -92 -1115 -80 -739
rect -138 -1127 -80 -1115
rect 80 -739 138 -727
rect 80 -1115 92 -739
rect 126 -1115 138 -739
rect 80 -1127 138 -1115
<< mvndiffc >>
rect -126 739 -92 1115
rect 92 739 126 1115
rect -126 121 -92 497
rect 92 121 126 497
rect -126 -497 -92 -121
rect 92 -497 126 -121
rect -126 -1115 -92 -739
rect 92 -1115 126 -739
<< mvpsubdiff >>
rect -272 1337 272 1349
rect -272 1303 -164 1337
rect 164 1303 272 1337
rect -272 1291 272 1303
rect -272 1241 -214 1291
rect -272 -1241 -260 1241
rect -226 -1241 -214 1241
rect 214 1241 272 1291
rect -272 -1291 -214 -1241
rect 214 -1241 226 1241
rect 260 -1241 272 1241
rect 214 -1291 272 -1241
rect -272 -1303 272 -1291
rect -272 -1337 -164 -1303
rect 164 -1337 272 -1303
rect -272 -1349 272 -1337
<< mvpsubdiffcont >>
rect -164 1303 164 1337
rect -260 -1241 -226 1241
rect 226 -1241 260 1241
rect -164 -1337 164 -1303
<< poly >>
rect -80 1199 80 1215
rect -80 1165 -64 1199
rect 64 1165 80 1199
rect -80 1127 80 1165
rect -80 689 80 727
rect -80 655 -64 689
rect 64 655 80 689
rect -80 639 80 655
rect -80 581 80 597
rect -80 547 -64 581
rect 64 547 80 581
rect -80 509 80 547
rect -80 71 80 109
rect -80 37 -64 71
rect 64 37 80 71
rect -80 21 80 37
rect -80 -37 80 -21
rect -80 -71 -64 -37
rect 64 -71 80 -37
rect -80 -109 80 -71
rect -80 -547 80 -509
rect -80 -581 -64 -547
rect 64 -581 80 -547
rect -80 -597 80 -581
rect -80 -655 80 -639
rect -80 -689 -64 -655
rect 64 -689 80 -655
rect -80 -727 80 -689
rect -80 -1165 80 -1127
rect -80 -1199 -64 -1165
rect 64 -1199 80 -1165
rect -80 -1215 80 -1199
<< polycont >>
rect -64 1165 64 1199
rect -64 655 64 689
rect -64 547 64 581
rect -64 37 64 71
rect -64 -71 64 -37
rect -64 -581 64 -547
rect -64 -689 64 -655
rect -64 -1199 64 -1165
<< locali >>
rect -260 1303 -164 1337
rect 164 1303 260 1337
rect -260 1241 -226 1303
rect 226 1241 260 1303
rect -80 1165 -64 1199
rect 64 1165 80 1199
rect -126 1115 -92 1131
rect -126 723 -92 739
rect 92 1115 126 1131
rect 92 723 126 739
rect -80 655 -64 689
rect 64 655 80 689
rect -80 547 -64 581
rect 64 547 80 581
rect -126 497 -92 513
rect -126 105 -92 121
rect 92 497 126 513
rect 92 105 126 121
rect -80 37 -64 71
rect 64 37 80 71
rect -80 -71 -64 -37
rect 64 -71 80 -37
rect -126 -121 -92 -105
rect -126 -513 -92 -497
rect 92 -121 126 -105
rect 92 -513 126 -497
rect -80 -581 -64 -547
rect 64 -581 80 -547
rect -80 -689 -64 -655
rect 64 -689 80 -655
rect -126 -739 -92 -723
rect -126 -1131 -92 -1115
rect 92 -739 126 -723
rect 92 -1131 126 -1115
rect -80 -1199 -64 -1165
rect 64 -1199 80 -1165
rect -260 -1303 -226 -1241
rect 226 -1303 260 -1241
rect -260 -1337 -164 -1303
rect 164 -1337 260 -1303
<< viali >>
rect -64 1165 64 1199
rect -126 739 -92 1115
rect 92 739 126 1115
rect -64 655 64 689
rect -64 547 64 581
rect -126 121 -92 497
rect 92 121 126 497
rect -64 37 64 71
rect -64 -71 64 -37
rect -126 -497 -92 -121
rect 92 -497 126 -121
rect -64 -581 64 -547
rect -64 -689 64 -655
rect -126 -1115 -92 -739
rect 92 -1115 126 -739
rect -64 -1199 64 -1165
<< metal1 >>
rect -76 1199 76 1205
rect -76 1165 -64 1199
rect 64 1165 76 1199
rect -76 1159 76 1165
rect -132 1115 -86 1127
rect -132 739 -126 1115
rect -92 739 -86 1115
rect -132 727 -86 739
rect 86 1115 132 1127
rect 86 739 92 1115
rect 126 739 132 1115
rect 86 727 132 739
rect -76 689 76 695
rect -76 655 -64 689
rect 64 655 76 689
rect -76 649 76 655
rect -76 581 76 587
rect -76 547 -64 581
rect 64 547 76 581
rect -76 541 76 547
rect -132 497 -86 509
rect -132 121 -126 497
rect -92 121 -86 497
rect -132 109 -86 121
rect 86 497 132 509
rect 86 121 92 497
rect 126 121 132 497
rect 86 109 132 121
rect -76 71 76 77
rect -76 37 -64 71
rect 64 37 76 71
rect -76 31 76 37
rect -76 -37 76 -31
rect -76 -71 -64 -37
rect 64 -71 76 -37
rect -76 -77 76 -71
rect -132 -121 -86 -109
rect -132 -497 -126 -121
rect -92 -497 -86 -121
rect -132 -509 -86 -497
rect 86 -121 132 -109
rect 86 -497 92 -121
rect 126 -497 132 -121
rect 86 -509 132 -497
rect -76 -547 76 -541
rect -76 -581 -64 -547
rect 64 -581 76 -547
rect -76 -587 76 -581
rect -76 -655 76 -649
rect -76 -689 -64 -655
rect 64 -689 76 -655
rect -76 -695 76 -689
rect -132 -739 -86 -727
rect -132 -1115 -126 -739
rect -92 -1115 -86 -739
rect -132 -1127 -86 -1115
rect 86 -739 132 -727
rect 86 -1115 92 -739
rect 126 -1115 132 -739
rect 86 -1127 132 -1115
rect -76 -1165 76 -1159
rect -76 -1199 -64 -1165
rect 64 -1199 76 -1165
rect -76 -1205 76 -1199
<< properties >>
string FIXED_BBOX -243 -1320 243 1320
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2.0 l 0.8 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
