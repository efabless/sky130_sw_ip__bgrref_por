magic
tech sky130A
magscale 1 2
timestamp 1717527227
<< metal4 >>
rect -1949 1639 1949 1680
rect -1949 -1639 1693 1639
rect 1929 -1639 1949 1639
rect -1949 -1680 1949 -1639
<< via4 >>
rect 1693 -1639 1929 1639
<< mimcap2 >>
rect -1869 1560 1331 1600
rect -1869 -1560 -1829 1560
rect 1291 -1560 1331 1560
rect -1869 -1600 1331 -1560
<< mimcap2contact >>
rect -1829 -1560 1291 1560
<< metal5 >>
rect 1651 1639 1971 1681
rect -1853 1560 1315 1584
rect -1853 -1560 -1829 1560
rect 1291 -1560 1315 1560
rect -1853 -1584 1315 -1560
rect 1651 -1639 1693 1639
rect 1929 -1639 1971 1639
rect 1651 -1681 1971 -1639
<< properties >>
string FIXED_BBOX -1949 -1680 1411 1680
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 16.0 l 16.0 val 524.159 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
