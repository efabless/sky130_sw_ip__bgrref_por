magic
tech sky130A
magscale 1 2
timestamp 1717527227
<< error_p >>
rect -88 138 -30 144
rect 30 138 88 144
rect -88 104 -76 138
rect 30 104 42 138
rect -88 98 -30 104
rect 30 98 88 104
rect -88 -104 -30 -98
rect 30 -104 88 -98
rect -88 -138 -76 -104
rect 30 -138 42 -104
rect -88 -144 -30 -138
rect 30 -144 88 -138
<< pwell >>
rect -285 -260 285 260
<< nmos >>
rect -89 -50 -29 50
rect 29 -50 89 50
<< ndiff >>
rect -147 38 -89 50
rect -147 -38 -135 38
rect -101 -38 -89 38
rect -147 -50 -89 -38
rect -29 38 29 50
rect -29 -38 -17 38
rect 17 -38 29 38
rect -29 -50 29 -38
rect 89 38 147 50
rect 89 -38 101 38
rect 135 -38 147 38
rect 89 -50 147 -38
<< ndiffc >>
rect -135 -38 -101 38
rect -17 -38 17 38
rect 101 -38 135 38
<< psubdiff >>
rect -249 190 -153 224
rect 153 190 249 224
rect -249 128 -215 190
rect 215 128 249 190
rect -249 -190 -215 -128
rect 215 -190 249 -128
rect -249 -224 -153 -190
rect 153 -224 249 -190
<< psubdiffcont >>
rect -153 190 153 224
rect -249 -128 -215 128
rect 215 -128 249 128
rect -153 -224 153 -190
<< poly >>
rect -92 138 -26 154
rect -92 104 -76 138
rect -42 104 -26 138
rect -92 88 -26 104
rect 26 138 92 154
rect 26 104 42 138
rect 76 104 92 138
rect 26 88 92 104
rect -89 50 -29 88
rect 29 50 89 88
rect -89 -88 -29 -50
rect 29 -88 89 -50
rect -92 -104 -26 -88
rect -92 -138 -76 -104
rect -42 -138 -26 -104
rect -92 -154 -26 -138
rect 26 -104 92 -88
rect 26 -138 42 -104
rect 76 -138 92 -104
rect 26 -154 92 -138
<< polycont >>
rect -76 104 -42 138
rect 42 104 76 138
rect -76 -138 -42 -104
rect 42 -138 76 -104
<< locali >>
rect -249 190 -153 224
rect 153 190 249 224
rect -249 128 -215 190
rect -92 104 -76 138
rect -42 104 -26 138
rect 26 104 42 138
rect 76 104 92 138
rect 215 128 249 190
rect -135 38 -101 54
rect -135 -54 -101 -38
rect -17 38 17 54
rect -17 -54 17 -38
rect 101 38 135 54
rect 101 -54 135 -38
rect -249 -190 -215 -128
rect -92 -138 -76 -104
rect -42 -138 -26 -104
rect 26 -138 42 -104
rect 76 -138 92 -104
rect 215 -190 249 -128
rect -249 -224 -153 -190
rect 153 -224 249 -190
<< viali >>
rect -76 104 -42 138
rect 42 104 76 138
rect -135 -38 -101 38
rect -17 -38 17 38
rect 101 -38 135 38
rect -76 -138 -42 -104
rect 42 -138 76 -104
<< metal1 >>
rect -88 138 -30 144
rect -88 104 -76 138
rect -42 104 -30 138
rect -88 98 -30 104
rect 30 138 88 144
rect 30 104 42 138
rect 76 104 88 138
rect 30 98 88 104
rect -141 38 -95 50
rect -141 -38 -135 38
rect -101 -38 -95 38
rect -141 -50 -95 -38
rect -23 38 23 50
rect -23 -38 -17 38
rect 17 -38 23 38
rect -23 -50 23 -38
rect 95 38 141 50
rect 95 -38 101 38
rect 135 -38 141 38
rect 95 -50 141 -38
rect -88 -104 -30 -98
rect -88 -138 -76 -104
rect -42 -138 -30 -104
rect -88 -144 -30 -138
rect 30 -104 88 -98
rect 30 -138 42 -104
rect 76 -138 88 -104
rect 30 -144 88 -138
<< properties >>
string FIXED_BBOX -232 -207 232 207
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.3 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
