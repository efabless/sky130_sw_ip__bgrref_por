magic
tech sky130A
magscale 1 2
timestamp 1717527227
<< nwell >>
rect 33421 -285686 33423 -285354
<< locali >>
rect 33368 -285226 33451 -285225
rect 33368 -285246 36265 -285226
rect 33368 -285285 33432 -285246
rect 36173 -285285 36265 -285246
rect 33368 -285320 36265 -285285
rect 33368 -285354 33451 -285320
rect 33368 -285686 33389 -285354
rect 33423 -285686 33451 -285354
rect 33368 -285710 33451 -285686
rect 36185 -285347 36265 -285320
rect 36185 -285850 36208 -285347
rect 36242 -285850 36265 -285347
rect 36185 -285895 36265 -285850
rect 36194 -286070 36258 -286034
rect 33372 -286251 33440 -286226
rect 33372 -286411 33386 -286251
rect 33421 -286411 33440 -286251
rect 33372 -286433 33440 -286411
rect 36194 -286411 36208 -286070
rect 36243 -286411 36258 -286070
rect 36194 -286433 36258 -286411
rect 33372 -286452 36258 -286433
rect 33372 -286491 33447 -286452
rect 36188 -286491 36258 -286452
rect 33372 -286515 36258 -286491
<< viali >>
rect 33432 -285285 36173 -285246
rect 33389 -285686 33423 -285354
rect 36208 -285850 36242 -285347
rect 33386 -286411 33421 -286251
rect 36208 -286411 36243 -286070
rect 33447 -286491 36188 -286452
<< metal1 >>
rect 33368 -285226 33451 -285225
rect 33368 -285241 36265 -285226
rect 33368 -285246 33440 -285241
rect 33368 -285285 33432 -285246
rect 33368 -285304 33440 -285285
rect 36182 -285304 36265 -285241
rect 33368 -285320 36265 -285304
rect 33368 -285354 33451 -285320
rect 33368 -285686 33389 -285354
rect 33423 -285686 33451 -285354
rect 33368 -285710 33451 -285686
rect 36185 -285347 36265 -285320
rect 33417 -285810 33524 -285764
rect 33417 -285917 33463 -285810
rect 33354 -286009 33463 -285917
rect 33417 -286140 33463 -286009
rect 33417 -286186 33522 -286140
rect 33614 -286185 33654 -285764
rect 33806 -286186 33846 -285764
rect 34574 -285940 34614 -285763
rect 36185 -285850 36208 -285347
rect 36242 -285850 36265 -285347
rect 36185 -285895 36265 -285850
rect 34506 -285992 34614 -285940
rect 34574 -286186 34614 -285992
rect 36194 -286070 36258 -286034
rect 33372 -286251 33440 -286226
rect 33372 -286411 33386 -286251
rect 33421 -286411 33440 -286251
rect 33372 -286433 33440 -286411
rect 36194 -286411 36208 -286070
rect 36243 -286411 36258 -286070
rect 36194 -286433 36258 -286411
rect 33372 -286441 36258 -286433
rect 33372 -286452 33449 -286441
rect 33372 -286491 33447 -286452
rect 33372 -286504 33449 -286491
rect 36191 -286504 36258 -286441
rect 33372 -286515 36258 -286504
<< via1 >>
rect 33440 -285246 36182 -285241
rect 33440 -285285 36173 -285246
rect 36173 -285285 36182 -285246
rect 33440 -285304 36182 -285285
rect 33449 -286452 36191 -286441
rect 33449 -286491 36188 -286452
rect 36188 -286491 36191 -286452
rect 33449 -286504 36191 -286491
<< metal2 >>
rect 33352 -285241 36280 -285202
rect 33352 -285304 33440 -285241
rect 36182 -285304 36280 -285241
rect 33352 -285357 36280 -285304
rect 33489 -286220 33553 -285387
rect 33585 -285392 33649 -285357
rect 33585 -285598 33649 -285514
rect 33681 -286220 33745 -285389
rect 33777 -285392 33841 -285357
rect 33777 -285598 33841 -285514
rect 33873 -285917 33937 -285389
rect 33969 -285392 34033 -285357
rect 33969 -285598 34033 -285514
rect 34065 -285917 34129 -285389
rect 34161 -285392 34225 -285357
rect 34161 -285598 34225 -285514
rect 34257 -285917 34321 -285389
rect 34353 -285392 34417 -285357
rect 34353 -285598 34417 -285514
rect 34449 -285917 34513 -285389
rect 34545 -285392 34609 -285357
rect 34545 -285598 34609 -285514
rect 33873 -286004 34513 -285917
rect 33873 -286220 33937 -286004
rect 34065 -286220 34129 -286004
rect 34257 -286220 34321 -286004
rect 34449 -286220 34513 -286004
rect 34641 -285917 34705 -285389
rect 34737 -285392 34801 -285357
rect 34737 -285598 34801 -285514
rect 34833 -285917 34897 -285389
rect 34929 -285392 34993 -285357
rect 34929 -285598 34993 -285514
rect 35025 -285917 35089 -285389
rect 35121 -285392 35185 -285357
rect 35121 -285598 35185 -285514
rect 35217 -285917 35281 -285389
rect 35313 -285392 35377 -285357
rect 35313 -285598 35377 -285514
rect 35409 -285917 35473 -285389
rect 35505 -285392 35569 -285357
rect 35505 -285598 35569 -285514
rect 35601 -285917 35665 -285389
rect 35697 -285392 35761 -285357
rect 35697 -285598 35761 -285514
rect 35793 -285917 35857 -285389
rect 35889 -285392 35953 -285357
rect 35889 -285598 35953 -285514
rect 35985 -285912 36049 -285389
rect 36081 -285392 36145 -285357
rect 36081 -285598 36145 -285514
rect 35985 -285917 36281 -285912
rect 34641 -286004 36281 -285917
rect 34641 -286220 34705 -286004
rect 34833 -286220 34897 -286004
rect 35025 -286220 35089 -286004
rect 35217 -286220 35281 -286004
rect 35409 -286220 35473 -286004
rect 35601 -286220 35665 -286004
rect 35793 -286220 35857 -286004
rect 35985 -286019 36281 -286004
rect 35985 -286220 36049 -286019
rect 33585 -286374 33649 -286342
rect 33777 -286374 33841 -286342
rect 33969 -286374 34033 -286342
rect 34161 -286374 34225 -286342
rect 34353 -286374 34417 -286342
rect 34545 -286374 34609 -286342
rect 34737 -286374 34801 -286342
rect 34929 -286374 34993 -286342
rect 35121 -286374 35185 -286342
rect 35313 -286374 35377 -286342
rect 35505 -286374 35569 -286342
rect 35697 -286374 35761 -286342
rect 35889 -286374 35953 -286342
rect 36081 -286374 36145 -286342
rect 33355 -286441 36280 -286374
rect 33355 -286504 33449 -286441
rect 36191 -286504 36280 -286441
rect 33355 -286527 36280 -286504
use por_via_2cut  por_via_2cut_0
timestamp 1717527227
transform 0 1 42573 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_1
timestamp 1717527227
transform 0 1 41421 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_2
timestamp 1717527227
transform 0 1 41421 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_3
timestamp 1717527227
transform 0 1 41613 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_4
timestamp 1717527227
transform 0 1 41517 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_5
timestamp 1717527227
transform 0 1 41709 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_6
timestamp 1717527227
transform 0 1 41805 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_7
timestamp 1717527227
transform 0 1 41901 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_8
timestamp 1717527227
transform 0 1 41997 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_9
timestamp 1717527227
transform 0 1 42093 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_10
timestamp 1717527227
transform 0 1 42189 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_11
timestamp 1717527227
transform 0 1 42285 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_12
timestamp 1717527227
transform 0 1 42381 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_13
timestamp 1717527227
transform 0 1 42477 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_14
timestamp 1717527227
transform 0 1 42861 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_15
timestamp 1717527227
transform 0 1 42669 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_16
timestamp 1717527227
transform 0 1 42765 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_17
timestamp 1717527227
transform 0 1 43053 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_18
timestamp 1717527227
transform 0 1 42957 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_19
timestamp 1717527227
transform 0 1 43341 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_20
timestamp 1717527227
transform 0 1 43149 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_21
timestamp 1717527227
transform 0 1 43245 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_22
timestamp 1717527227
transform 0 1 43629 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_23
timestamp 1717527227
transform 0 1 43437 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_24
timestamp 1717527227
transform 0 1 43533 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_25
timestamp 1717527227
transform 0 1 43917 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_26
timestamp 1717527227
transform 0 1 43725 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_27
timestamp 1717527227
transform 0 1 43821 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_28
timestamp 1717527227
transform 0 1 44013 -1 0 -270126
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_29
timestamp 1717527227
transform 0 1 42381 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_30
timestamp 1717527227
transform 0 1 42381 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_31
timestamp 1717527227
transform -1 0 49714 0 -1 -293867
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_32
timestamp 1717527227
transform 0 1 41421 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_33
timestamp 1717527227
transform 0 1 41517 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_34
timestamp 1717527227
transform 0 1 41517 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_35
timestamp 1717527227
transform 0 1 41613 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_36
timestamp 1717527227
transform 0 1 41613 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_37
timestamp 1717527227
transform 0 1 41709 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_38
timestamp 1717527227
transform 0 1 41709 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_39
timestamp 1717527227
transform 0 1 41805 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_40
timestamp 1717527227
transform 0 1 41805 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_41
timestamp 1717527227
transform 0 1 41901 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_42
timestamp 1717527227
transform 0 1 41901 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_43
timestamp 1717527227
transform 0 1 41997 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_44
timestamp 1717527227
transform 0 1 41997 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_45
timestamp 1717527227
transform 0 1 42093 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_46
timestamp 1717527227
transform 0 1 42093 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_47
timestamp 1717527227
transform 0 1 42189 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_48
timestamp 1717527227
transform 0 1 42189 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_49
timestamp 1717527227
transform 0 1 42285 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_50
timestamp 1717527227
transform 0 1 42285 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_51
timestamp 1717527227
transform 0 1 42669 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_52
timestamp 1717527227
transform 0 1 42669 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_53
timestamp 1717527227
transform 0 1 42477 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_54
timestamp 1717527227
transform 0 1 42477 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_55
timestamp 1717527227
transform 0 1 42573 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_56
timestamp 1717527227
transform 0 1 42573 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_57
timestamp 1717527227
transform 0 1 42957 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_58
timestamp 1717527227
transform 0 1 42957 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_59
timestamp 1717527227
transform 0 1 42765 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_60
timestamp 1717527227
transform 0 1 42765 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_61
timestamp 1717527227
transform 0 1 42861 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_62
timestamp 1717527227
transform 0 1 42861 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_63
timestamp 1717527227
transform 0 1 43245 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_64
timestamp 1717527227
transform 0 1 43245 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_65
timestamp 1717527227
transform 0 1 43053 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_66
timestamp 1717527227
transform 0 1 43053 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_67
timestamp 1717527227
transform 0 1 43149 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_68
timestamp 1717527227
transform 0 1 43149 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_69
timestamp 1717527227
transform 0 1 43629 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_70
timestamp 1717527227
transform 0 1 43629 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_71
timestamp 1717527227
transform 0 1 43341 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_72
timestamp 1717527227
transform 0 1 43341 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_73
timestamp 1717527227
transform 0 1 43437 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_74
timestamp 1717527227
transform 0 1 43437 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_75
timestamp 1717527227
transform 0 1 43533 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_76
timestamp 1717527227
transform 0 1 43533 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_77
timestamp 1717527227
transform 0 1 43917 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_78
timestamp 1717527227
transform 0 1 43917 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_79
timestamp 1717527227
transform 0 1 43725 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_80
timestamp 1717527227
transform 0 1 43725 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_81
timestamp 1717527227
transform 0 1 43821 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_82
timestamp 1717527227
transform 0 1 43821 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_83
timestamp 1717527227
transform 0 1 44013 -1 0 -269504
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_84
timestamp 1717527227
transform 0 1 44013 -1 0 -269298
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_85
timestamp 1717527227
transform -1 0 49905 0 -1 -293868
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_86
timestamp 1717527227
transform -1 0 50594 0 -1 -293866
box 16088 -7932 16222 -7868
use sky130_fd_pr__nfet_01v8_PR763Z  XM53
timestamp 1717527227
transform 1 0 34817 0 1 -286268
box -1463 -260 1463 260
use sky130_fd_pr__pfet_01v8_DD63S8  XM54
timestamp 1717527227
transform 1 0 34819 0 1 -285521
box -1463 -397 1463 297
<< end >>
