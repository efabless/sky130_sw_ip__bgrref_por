magic
tech sky130A
magscale 1 2
timestamp 1717527227
<< metal4 >>
rect -21290 3439 -17392 3480
rect -21290 161 -17648 3439
rect -17412 161 -17392 3439
rect -21290 120 -17392 161
rect -16992 3439 -13094 3480
rect -16992 161 -13350 3439
rect -13114 161 -13094 3439
rect -16992 120 -13094 161
rect -12694 3439 -8796 3480
rect -12694 161 -9052 3439
rect -8816 161 -8796 3439
rect -12694 120 -8796 161
rect -8396 3439 -4498 3480
rect -8396 161 -4754 3439
rect -4518 161 -4498 3439
rect -8396 120 -4498 161
rect -4098 3439 -200 3480
rect -4098 161 -456 3439
rect -220 161 -200 3439
rect -4098 120 -200 161
rect 200 3439 4098 3480
rect 200 161 3842 3439
rect 4078 161 4098 3439
rect 200 120 4098 161
rect 4498 3439 8396 3480
rect 4498 161 8140 3439
rect 8376 161 8396 3439
rect 4498 120 8396 161
rect 8796 3439 12694 3480
rect 8796 161 12438 3439
rect 12674 161 12694 3439
rect 8796 120 12694 161
rect 13094 3439 16992 3480
rect 13094 161 16736 3439
rect 16972 161 16992 3439
rect 13094 120 16992 161
rect 17392 3439 21290 3480
rect 17392 161 21034 3439
rect 21270 161 21290 3439
rect 17392 120 21290 161
rect -21290 -161 -17392 -120
rect -21290 -3439 -17648 -161
rect -17412 -3439 -17392 -161
rect -21290 -3480 -17392 -3439
rect -16992 -161 -13094 -120
rect -16992 -3439 -13350 -161
rect -13114 -3439 -13094 -161
rect -16992 -3480 -13094 -3439
rect -12694 -161 -8796 -120
rect -12694 -3439 -9052 -161
rect -8816 -3439 -8796 -161
rect -12694 -3480 -8796 -3439
rect -8396 -161 -4498 -120
rect -8396 -3439 -4754 -161
rect -4518 -3439 -4498 -161
rect -8396 -3480 -4498 -3439
rect -4098 -161 -200 -120
rect -4098 -3439 -456 -161
rect -220 -3439 -200 -161
rect -4098 -3480 -200 -3439
rect 200 -161 4098 -120
rect 200 -3439 3842 -161
rect 4078 -3439 4098 -161
rect 200 -3480 4098 -3439
rect 4498 -161 8396 -120
rect 4498 -3439 8140 -161
rect 8376 -3439 8396 -161
rect 4498 -3480 8396 -3439
rect 8796 -161 12694 -120
rect 8796 -3439 12438 -161
rect 12674 -3439 12694 -161
rect 8796 -3480 12694 -3439
rect 13094 -161 16992 -120
rect 13094 -3439 16736 -161
rect 16972 -3439 16992 -161
rect 13094 -3480 16992 -3439
rect 17392 -161 21290 -120
rect 17392 -3439 21034 -161
rect 21270 -3439 21290 -161
rect 17392 -3480 21290 -3439
<< via4 >>
rect -17648 161 -17412 3439
rect -13350 161 -13114 3439
rect -9052 161 -8816 3439
rect -4754 161 -4518 3439
rect -456 161 -220 3439
rect 3842 161 4078 3439
rect 8140 161 8376 3439
rect 12438 161 12674 3439
rect 16736 161 16972 3439
rect 21034 161 21270 3439
rect -17648 -3439 -17412 -161
rect -13350 -3439 -13114 -161
rect -9052 -3439 -8816 -161
rect -4754 -3439 -4518 -161
rect -456 -3439 -220 -161
rect 3842 -3439 4078 -161
rect 8140 -3439 8376 -161
rect 12438 -3439 12674 -161
rect 16736 -3439 16972 -161
rect 21034 -3439 21270 -161
<< mimcap2 >>
rect -21210 3360 -18010 3400
rect -21210 240 -21170 3360
rect -18050 240 -18010 3360
rect -21210 200 -18010 240
rect -16912 3360 -13712 3400
rect -16912 240 -16872 3360
rect -13752 240 -13712 3360
rect -16912 200 -13712 240
rect -12614 3360 -9414 3400
rect -12614 240 -12574 3360
rect -9454 240 -9414 3360
rect -12614 200 -9414 240
rect -8316 3360 -5116 3400
rect -8316 240 -8276 3360
rect -5156 240 -5116 3360
rect -8316 200 -5116 240
rect -4018 3360 -818 3400
rect -4018 240 -3978 3360
rect -858 240 -818 3360
rect -4018 200 -818 240
rect 280 3360 3480 3400
rect 280 240 320 3360
rect 3440 240 3480 3360
rect 280 200 3480 240
rect 4578 3360 7778 3400
rect 4578 240 4618 3360
rect 7738 240 7778 3360
rect 4578 200 7778 240
rect 8876 3360 12076 3400
rect 8876 240 8916 3360
rect 12036 240 12076 3360
rect 8876 200 12076 240
rect 13174 3360 16374 3400
rect 13174 240 13214 3360
rect 16334 240 16374 3360
rect 13174 200 16374 240
rect 17472 3360 20672 3400
rect 17472 240 17512 3360
rect 20632 240 20672 3360
rect 17472 200 20672 240
rect -21210 -240 -18010 -200
rect -21210 -3360 -21170 -240
rect -18050 -3360 -18010 -240
rect -21210 -3400 -18010 -3360
rect -16912 -240 -13712 -200
rect -16912 -3360 -16872 -240
rect -13752 -3360 -13712 -240
rect -16912 -3400 -13712 -3360
rect -12614 -240 -9414 -200
rect -12614 -3360 -12574 -240
rect -9454 -3360 -9414 -240
rect -12614 -3400 -9414 -3360
rect -8316 -240 -5116 -200
rect -8316 -3360 -8276 -240
rect -5156 -3360 -5116 -240
rect -8316 -3400 -5116 -3360
rect -4018 -240 -818 -200
rect -4018 -3360 -3978 -240
rect -858 -3360 -818 -240
rect -4018 -3400 -818 -3360
rect 280 -240 3480 -200
rect 280 -3360 320 -240
rect 3440 -3360 3480 -240
rect 280 -3400 3480 -3360
rect 4578 -240 7778 -200
rect 4578 -3360 4618 -240
rect 7738 -3360 7778 -240
rect 4578 -3400 7778 -3360
rect 8876 -240 12076 -200
rect 8876 -3360 8916 -240
rect 12036 -3360 12076 -240
rect 8876 -3400 12076 -3360
rect 13174 -240 16374 -200
rect 13174 -3360 13214 -240
rect 16334 -3360 16374 -240
rect 13174 -3400 16374 -3360
rect 17472 -240 20672 -200
rect 17472 -3360 17512 -240
rect 20632 -3360 20672 -240
rect 17472 -3400 20672 -3360
<< mimcap2contact >>
rect -21170 240 -18050 3360
rect -16872 240 -13752 3360
rect -12574 240 -9454 3360
rect -8276 240 -5156 3360
rect -3978 240 -858 3360
rect 320 240 3440 3360
rect 4618 240 7738 3360
rect 8916 240 12036 3360
rect 13214 240 16334 3360
rect 17512 240 20632 3360
rect -21170 -3360 -18050 -240
rect -16872 -3360 -13752 -240
rect -12574 -3360 -9454 -240
rect -8276 -3360 -5156 -240
rect -3978 -3360 -858 -240
rect 320 -3360 3440 -240
rect 4618 -3360 7738 -240
rect 8916 -3360 12036 -240
rect 13214 -3360 16334 -240
rect 17512 -3360 20632 -240
<< metal5 >>
rect -19770 3384 -19450 3600
rect -17690 3439 -17370 3600
rect -21194 3360 -18026 3384
rect -21194 240 -21170 3360
rect -18050 240 -18026 3360
rect -21194 216 -18026 240
rect -19770 -216 -19450 216
rect -17690 161 -17648 3439
rect -17412 161 -17370 3439
rect -15472 3384 -15152 3600
rect -13392 3439 -13072 3600
rect -16896 3360 -13728 3384
rect -16896 240 -16872 3360
rect -13752 240 -13728 3360
rect -16896 216 -13728 240
rect -17690 -161 -17370 161
rect -21194 -240 -18026 -216
rect -21194 -3360 -21170 -240
rect -18050 -3360 -18026 -240
rect -21194 -3384 -18026 -3360
rect -19770 -3600 -19450 -3384
rect -17690 -3439 -17648 -161
rect -17412 -3439 -17370 -161
rect -15472 -216 -15152 216
rect -13392 161 -13350 3439
rect -13114 161 -13072 3439
rect -11174 3384 -10854 3600
rect -9094 3439 -8774 3600
rect -12598 3360 -9430 3384
rect -12598 240 -12574 3360
rect -9454 240 -9430 3360
rect -12598 216 -9430 240
rect -13392 -161 -13072 161
rect -16896 -240 -13728 -216
rect -16896 -3360 -16872 -240
rect -13752 -3360 -13728 -240
rect -16896 -3384 -13728 -3360
rect -17690 -3600 -17370 -3439
rect -15472 -3600 -15152 -3384
rect -13392 -3439 -13350 -161
rect -13114 -3439 -13072 -161
rect -11174 -216 -10854 216
rect -9094 161 -9052 3439
rect -8816 161 -8774 3439
rect -6876 3384 -6556 3600
rect -4796 3439 -4476 3600
rect -8300 3360 -5132 3384
rect -8300 240 -8276 3360
rect -5156 240 -5132 3360
rect -8300 216 -5132 240
rect -9094 -161 -8774 161
rect -12598 -240 -9430 -216
rect -12598 -3360 -12574 -240
rect -9454 -3360 -9430 -240
rect -12598 -3384 -9430 -3360
rect -13392 -3600 -13072 -3439
rect -11174 -3600 -10854 -3384
rect -9094 -3439 -9052 -161
rect -8816 -3439 -8774 -161
rect -6876 -216 -6556 216
rect -4796 161 -4754 3439
rect -4518 161 -4476 3439
rect -2578 3384 -2258 3600
rect -498 3439 -178 3600
rect -4002 3360 -834 3384
rect -4002 240 -3978 3360
rect -858 240 -834 3360
rect -4002 216 -834 240
rect -4796 -161 -4476 161
rect -8300 -240 -5132 -216
rect -8300 -3360 -8276 -240
rect -5156 -3360 -5132 -240
rect -8300 -3384 -5132 -3360
rect -9094 -3600 -8774 -3439
rect -6876 -3600 -6556 -3384
rect -4796 -3439 -4754 -161
rect -4518 -3439 -4476 -161
rect -2578 -216 -2258 216
rect -498 161 -456 3439
rect -220 161 -178 3439
rect 1720 3384 2040 3600
rect 3800 3439 4120 3600
rect 296 3360 3464 3384
rect 296 240 320 3360
rect 3440 240 3464 3360
rect 296 216 3464 240
rect -498 -161 -178 161
rect -4002 -240 -834 -216
rect -4002 -3360 -3978 -240
rect -858 -3360 -834 -240
rect -4002 -3384 -834 -3360
rect -4796 -3600 -4476 -3439
rect -2578 -3600 -2258 -3384
rect -498 -3439 -456 -161
rect -220 -3439 -178 -161
rect 1720 -216 2040 216
rect 3800 161 3842 3439
rect 4078 161 4120 3439
rect 6018 3384 6338 3600
rect 8098 3439 8418 3600
rect 4594 3360 7762 3384
rect 4594 240 4618 3360
rect 7738 240 7762 3360
rect 4594 216 7762 240
rect 3800 -161 4120 161
rect 296 -240 3464 -216
rect 296 -3360 320 -240
rect 3440 -3360 3464 -240
rect 296 -3384 3464 -3360
rect -498 -3600 -178 -3439
rect 1720 -3600 2040 -3384
rect 3800 -3439 3842 -161
rect 4078 -3439 4120 -161
rect 6018 -216 6338 216
rect 8098 161 8140 3439
rect 8376 161 8418 3439
rect 10316 3384 10636 3600
rect 12396 3439 12716 3600
rect 8892 3360 12060 3384
rect 8892 240 8916 3360
rect 12036 240 12060 3360
rect 8892 216 12060 240
rect 8098 -161 8418 161
rect 4594 -240 7762 -216
rect 4594 -3360 4618 -240
rect 7738 -3360 7762 -240
rect 4594 -3384 7762 -3360
rect 3800 -3600 4120 -3439
rect 6018 -3600 6338 -3384
rect 8098 -3439 8140 -161
rect 8376 -3439 8418 -161
rect 10316 -216 10636 216
rect 12396 161 12438 3439
rect 12674 161 12716 3439
rect 14614 3384 14934 3600
rect 16694 3439 17014 3600
rect 13190 3360 16358 3384
rect 13190 240 13214 3360
rect 16334 240 16358 3360
rect 13190 216 16358 240
rect 12396 -161 12716 161
rect 8892 -240 12060 -216
rect 8892 -3360 8916 -240
rect 12036 -3360 12060 -240
rect 8892 -3384 12060 -3360
rect 8098 -3600 8418 -3439
rect 10316 -3600 10636 -3384
rect 12396 -3439 12438 -161
rect 12674 -3439 12716 -161
rect 14614 -216 14934 216
rect 16694 161 16736 3439
rect 16972 161 17014 3439
rect 18912 3384 19232 3600
rect 20992 3439 21312 3600
rect 17488 3360 20656 3384
rect 17488 240 17512 3360
rect 20632 240 20656 3360
rect 17488 216 20656 240
rect 16694 -161 17014 161
rect 13190 -240 16358 -216
rect 13190 -3360 13214 -240
rect 16334 -3360 16358 -240
rect 13190 -3384 16358 -3360
rect 12396 -3600 12716 -3439
rect 14614 -3600 14934 -3384
rect 16694 -3439 16736 -161
rect 16972 -3439 17014 -161
rect 18912 -216 19232 216
rect 20992 161 21034 3439
rect 21270 161 21312 3439
rect 20992 -161 21312 161
rect 17488 -240 20656 -216
rect 17488 -3360 17512 -240
rect 20632 -3360 20656 -240
rect 17488 -3384 20656 -3360
rect 16694 -3600 17014 -3439
rect 18912 -3600 19232 -3384
rect 20992 -3439 21034 -161
rect 21270 -3439 21312 -161
rect 20992 -3600 21312 -3439
<< properties >>
string FIXED_BBOX 17392 120 20752 3480
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 16.0 l 16.0 val 524.159 carea 2.00 cperi 0.19 nx 10 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
