magic
tech sky130A
magscale 1 2
timestamp 1717527227
<< error_p >>
rect -1295 -249 -1237 -243
rect -1295 -283 -1283 -249
rect -1295 -289 -1237 -283
<< nwell >>
rect -1463 -397 1463 297
<< pmos >>
rect -1263 18 -1233 158
rect -1167 18 -1137 158
rect -1071 18 -1041 158
rect -975 18 -945 158
rect -879 18 -849 158
rect -783 18 -753 158
rect -687 18 -657 158
rect -591 18 -561 158
rect -495 18 -465 158
rect -399 18 -369 158
rect -303 18 -273 158
rect -207 18 -177 158
rect -111 18 -81 158
rect -15 18 15 158
rect 81 18 111 158
rect 177 18 207 158
rect 273 18 303 158
rect 369 18 399 158
rect 465 18 495 158
rect 561 18 591 158
rect 657 18 687 158
rect 753 18 783 158
rect 849 18 879 158
rect 945 18 975 158
rect 1041 18 1071 158
rect 1137 18 1167 158
rect 1233 18 1263 158
rect -1263 -202 -1233 -62
rect -1167 -202 -1137 -62
rect -1071 -202 -1041 -62
rect -975 -202 -945 -62
rect -879 -202 -849 -62
rect -783 -202 -753 -62
rect -687 -202 -657 -62
rect -591 -202 -561 -62
rect -495 -202 -465 -62
rect -399 -202 -369 -62
rect -303 -202 -273 -62
rect -207 -202 -177 -62
rect -111 -202 -81 -62
rect -15 -202 15 -62
rect 81 -202 111 -62
rect 177 -202 207 -62
rect 273 -202 303 -62
rect 369 -202 399 -62
rect 465 -202 495 -62
rect 561 -202 591 -62
rect 657 -202 687 -62
rect 753 -202 783 -62
rect 849 -202 879 -62
rect 945 -202 975 -62
rect 1041 -202 1071 -62
rect 1137 -202 1167 -62
rect 1233 -202 1263 -62
<< pdiff >>
rect -1325 146 -1263 158
rect -1325 30 -1313 146
rect -1279 30 -1263 146
rect -1325 18 -1263 30
rect -1233 146 -1167 158
rect -1233 30 -1217 146
rect -1183 30 -1167 146
rect -1233 18 -1167 30
rect -1137 146 -1071 158
rect -1137 30 -1121 146
rect -1087 30 -1071 146
rect -1137 18 -1071 30
rect -1041 146 -975 158
rect -1041 30 -1025 146
rect -991 30 -975 146
rect -1041 18 -975 30
rect -945 146 -879 158
rect -945 30 -929 146
rect -895 30 -879 146
rect -945 18 -879 30
rect -849 146 -783 158
rect -849 30 -833 146
rect -799 30 -783 146
rect -849 18 -783 30
rect -753 146 -687 158
rect -753 30 -737 146
rect -703 30 -687 146
rect -753 18 -687 30
rect -657 146 -591 158
rect -657 30 -641 146
rect -607 30 -591 146
rect -657 18 -591 30
rect -561 146 -495 158
rect -561 30 -545 146
rect -511 30 -495 146
rect -561 18 -495 30
rect -465 146 -399 158
rect -465 30 -449 146
rect -415 30 -399 146
rect -465 18 -399 30
rect -369 146 -303 158
rect -369 30 -353 146
rect -319 30 -303 146
rect -369 18 -303 30
rect -273 146 -207 158
rect -273 30 -257 146
rect -223 30 -207 146
rect -273 18 -207 30
rect -177 146 -111 158
rect -177 30 -161 146
rect -127 30 -111 146
rect -177 18 -111 30
rect -81 146 -15 158
rect -81 30 -65 146
rect -31 30 -15 146
rect -81 18 -15 30
rect 15 146 81 158
rect 15 30 31 146
rect 65 30 81 146
rect 15 18 81 30
rect 111 146 177 158
rect 111 30 127 146
rect 161 30 177 146
rect 111 18 177 30
rect 207 146 273 158
rect 207 30 223 146
rect 257 30 273 146
rect 207 18 273 30
rect 303 146 369 158
rect 303 30 319 146
rect 353 30 369 146
rect 303 18 369 30
rect 399 146 465 158
rect 399 30 415 146
rect 449 30 465 146
rect 399 18 465 30
rect 495 146 561 158
rect 495 30 511 146
rect 545 30 561 146
rect 495 18 561 30
rect 591 146 657 158
rect 591 30 607 146
rect 641 30 657 146
rect 591 18 657 30
rect 687 146 753 158
rect 687 30 703 146
rect 737 30 753 146
rect 687 18 753 30
rect 783 146 849 158
rect 783 30 799 146
rect 833 30 849 146
rect 783 18 849 30
rect 879 146 945 158
rect 879 30 895 146
rect 929 30 945 146
rect 879 18 945 30
rect 975 146 1041 158
rect 975 30 991 146
rect 1025 30 1041 146
rect 975 18 1041 30
rect 1071 146 1137 158
rect 1071 30 1087 146
rect 1121 30 1137 146
rect 1071 18 1137 30
rect 1167 146 1233 158
rect 1167 30 1183 146
rect 1217 30 1233 146
rect 1167 18 1233 30
rect 1263 146 1325 158
rect 1263 30 1279 146
rect 1313 30 1325 146
rect 1263 18 1325 30
rect -1325 -74 -1263 -62
rect -1325 -190 -1313 -74
rect -1279 -190 -1263 -74
rect -1325 -202 -1263 -190
rect -1233 -74 -1167 -62
rect -1233 -190 -1217 -74
rect -1183 -190 -1167 -74
rect -1233 -202 -1167 -190
rect -1137 -74 -1071 -62
rect -1137 -190 -1121 -74
rect -1087 -190 -1071 -74
rect -1137 -202 -1071 -190
rect -1041 -74 -975 -62
rect -1041 -190 -1025 -74
rect -991 -190 -975 -74
rect -1041 -202 -975 -190
rect -945 -74 -879 -62
rect -945 -190 -929 -74
rect -895 -190 -879 -74
rect -945 -202 -879 -190
rect -849 -74 -783 -62
rect -849 -190 -833 -74
rect -799 -190 -783 -74
rect -849 -202 -783 -190
rect -753 -74 -687 -62
rect -753 -190 -737 -74
rect -703 -190 -687 -74
rect -753 -202 -687 -190
rect -657 -74 -591 -62
rect -657 -190 -641 -74
rect -607 -190 -591 -74
rect -657 -202 -591 -190
rect -561 -74 -495 -62
rect -561 -190 -545 -74
rect -511 -190 -495 -74
rect -561 -202 -495 -190
rect -465 -74 -399 -62
rect -465 -190 -449 -74
rect -415 -190 -399 -74
rect -465 -202 -399 -190
rect -369 -74 -303 -62
rect -369 -190 -353 -74
rect -319 -190 -303 -74
rect -369 -202 -303 -190
rect -273 -74 -207 -62
rect -273 -190 -257 -74
rect -223 -190 -207 -74
rect -273 -202 -207 -190
rect -177 -74 -111 -62
rect -177 -190 -161 -74
rect -127 -190 -111 -74
rect -177 -202 -111 -190
rect -81 -74 -15 -62
rect -81 -190 -65 -74
rect -31 -190 -15 -74
rect -81 -202 -15 -190
rect 15 -74 81 -62
rect 15 -190 31 -74
rect 65 -190 81 -74
rect 15 -202 81 -190
rect 111 -74 177 -62
rect 111 -190 127 -74
rect 161 -190 177 -74
rect 111 -202 177 -190
rect 207 -74 273 -62
rect 207 -190 223 -74
rect 257 -190 273 -74
rect 207 -202 273 -190
rect 303 -74 369 -62
rect 303 -190 319 -74
rect 353 -190 369 -74
rect 303 -202 369 -190
rect 399 -74 465 -62
rect 399 -190 415 -74
rect 449 -190 465 -74
rect 399 -202 465 -190
rect 495 -74 561 -62
rect 495 -190 511 -74
rect 545 -190 561 -74
rect 495 -202 561 -190
rect 591 -74 657 -62
rect 591 -190 607 -74
rect 641 -190 657 -74
rect 591 -202 657 -190
rect 687 -74 753 -62
rect 687 -190 703 -74
rect 737 -190 753 -74
rect 687 -202 753 -190
rect 783 -74 849 -62
rect 783 -190 799 -74
rect 833 -190 849 -74
rect 783 -202 849 -190
rect 879 -74 945 -62
rect 879 -190 895 -74
rect 929 -190 945 -74
rect 879 -202 945 -190
rect 975 -74 1041 -62
rect 975 -190 991 -74
rect 1025 -190 1041 -74
rect 975 -202 1041 -190
rect 1071 -74 1137 -62
rect 1071 -190 1087 -74
rect 1121 -190 1137 -74
rect 1071 -202 1137 -190
rect 1167 -74 1233 -62
rect 1167 -190 1183 -74
rect 1217 -190 1233 -74
rect 1167 -202 1233 -190
rect 1263 -74 1325 -62
rect 1263 -190 1279 -74
rect 1313 -190 1325 -74
rect 1263 -202 1325 -190
<< pdiffc >>
rect -1313 30 -1279 146
rect -1217 30 -1183 146
rect -1121 30 -1087 146
rect -1025 30 -991 146
rect -929 30 -895 146
rect -833 30 -799 146
rect -737 30 -703 146
rect -641 30 -607 146
rect -545 30 -511 146
rect -449 30 -415 146
rect -353 30 -319 146
rect -257 30 -223 146
rect -161 30 -127 146
rect -65 30 -31 146
rect 31 30 65 146
rect 127 30 161 146
rect 223 30 257 146
rect 319 30 353 146
rect 415 30 449 146
rect 511 30 545 146
rect 607 30 641 146
rect 703 30 737 146
rect 799 30 833 146
rect 895 30 929 146
rect 991 30 1025 146
rect 1087 30 1121 146
rect 1183 30 1217 146
rect 1279 30 1313 146
rect -1313 -190 -1279 -74
rect -1217 -190 -1183 -74
rect -1121 -190 -1087 -74
rect -1025 -190 -991 -74
rect -929 -190 -895 -74
rect -833 -190 -799 -74
rect -737 -190 -703 -74
rect -641 -190 -607 -74
rect -545 -190 -511 -74
rect -449 -190 -415 -74
rect -353 -190 -319 -74
rect -257 -190 -223 -74
rect -161 -190 -127 -74
rect -65 -190 -31 -74
rect 31 -190 65 -74
rect 127 -190 161 -74
rect 223 -190 257 -74
rect 319 -190 353 -74
rect 415 -190 449 -74
rect 511 -190 545 -74
rect 607 -190 641 -74
rect 703 -190 737 -74
rect 799 -190 833 -74
rect 895 -190 929 -74
rect 991 -190 1025 -74
rect 1087 -190 1121 -74
rect 1183 -190 1217 -74
rect 1279 -190 1313 -74
<< nsubdiff >>
rect -1427 227 -1331 261
rect 1331 227 1427 261
rect -1427 165 -1393 227
rect 1393 165 1427 227
rect -1427 -327 -1393 -265
rect 1393 -327 1427 -265
rect -1427 -361 -1331 -327
rect 1331 -361 1427 -327
<< nsubdiffcont >>
rect -1331 227 1331 261
rect -1427 -265 -1393 165
rect 1393 -265 1427 165
rect -1331 -361 1331 -327
<< poly >>
rect -1263 158 -1233 189
rect -1167 158 -1137 189
rect -1071 158 -1041 189
rect -975 158 -945 189
rect -879 158 -849 189
rect -783 158 -753 189
rect -687 158 -657 189
rect -591 158 -561 189
rect -495 158 -465 189
rect -399 158 -369 189
rect -303 158 -273 189
rect -207 158 -177 189
rect -111 158 -81 189
rect -15 158 15 189
rect 81 158 111 189
rect 177 158 207 189
rect 273 158 303 189
rect 369 158 399 189
rect 465 158 495 189
rect 561 158 591 189
rect 657 158 687 189
rect 753 158 783 189
rect 849 158 879 189
rect 945 158 975 189
rect 1041 158 1071 189
rect 1137 158 1167 189
rect 1233 158 1263 189
rect -1263 -62 -1233 18
rect -1167 -62 -1137 18
rect -1071 -62 -1041 18
rect -975 -62 -945 18
rect -879 -62 -849 18
rect -783 -62 -753 18
rect -687 -62 -657 18
rect -591 -62 -561 18
rect -495 -62 -465 18
rect -399 -62 -369 18
rect -303 -62 -273 18
rect -207 -62 -177 18
rect -111 -62 -81 18
rect -15 -62 15 18
rect 81 -62 111 18
rect 177 -62 207 18
rect 273 -62 303 18
rect 369 -62 399 18
rect 465 -62 495 18
rect 561 -62 591 18
rect 657 -62 687 18
rect 753 -62 783 18
rect 849 -62 879 18
rect 945 -62 975 18
rect 1041 -62 1071 18
rect 1137 -62 1167 18
rect 1233 -62 1263 18
rect -1263 -233 -1233 -202
rect -1299 -249 -1233 -233
rect -1299 -283 -1283 -249
rect -1249 -283 -1233 -249
rect -1299 -299 -1233 -283
rect -1167 -233 -1137 -202
rect -1071 -233 -1041 -202
rect -1167 -249 -1041 -233
rect -1167 -283 -1151 -249
rect -1057 -283 -1041 -249
rect -1167 -299 -1041 -283
rect -975 -233 -945 -202
rect -879 -233 -849 -202
rect -783 -233 -753 -202
rect -687 -233 -657 -202
rect -591 -233 -561 -202
rect -495 -233 -465 -202
rect -399 -233 -369 -202
rect -303 -233 -273 -202
rect -975 -249 -273 -233
rect -975 -283 -959 -249
rect -289 -283 -273 -249
rect -975 -299 -273 -283
rect -207 -233 -177 -202
rect -111 -233 -81 -202
rect -15 -233 15 -202
rect 81 -233 111 -202
rect 177 -233 207 -202
rect 273 -233 303 -202
rect 369 -233 399 -202
rect 465 -233 495 -202
rect 561 -233 591 -202
rect 657 -233 687 -202
rect 753 -233 783 -202
rect 849 -233 879 -202
rect 945 -233 975 -202
rect 1041 -233 1071 -202
rect 1137 -233 1167 -202
rect 1233 -233 1263 -202
rect -207 -249 1263 -233
rect -207 -283 -191 -249
rect 1247 -283 1263 -249
rect -207 -299 1263 -283
<< polycont >>
rect -1283 -283 -1249 -249
rect -1151 -283 -1057 -249
rect -959 -283 -289 -249
rect -191 -283 1247 -249
<< locali >>
rect -1427 227 -1331 261
rect 1331 227 1427 261
rect -1427 165 -1393 227
rect 1393 165 1427 227
rect -1313 146 -1279 162
rect -1313 14 -1279 30
rect -1217 146 -1183 162
rect -1217 14 -1183 30
rect -1121 146 -1087 162
rect -1121 14 -1087 30
rect -1025 146 -991 162
rect -1025 14 -991 30
rect -929 146 -895 162
rect -929 14 -895 30
rect -833 146 -799 162
rect -833 14 -799 30
rect -737 146 -703 162
rect -737 14 -703 30
rect -641 146 -607 162
rect -641 14 -607 30
rect -545 146 -511 162
rect -545 14 -511 30
rect -449 146 -415 162
rect -449 14 -415 30
rect -353 146 -319 162
rect -353 14 -319 30
rect -257 146 -223 162
rect -257 14 -223 30
rect -161 146 -127 162
rect -161 14 -127 30
rect -65 146 -31 162
rect -65 14 -31 30
rect 31 146 65 162
rect 31 14 65 30
rect 127 146 161 162
rect 127 14 161 30
rect 223 146 257 162
rect 223 14 257 30
rect 319 146 353 162
rect 319 14 353 30
rect 415 146 449 162
rect 415 14 449 30
rect 511 146 545 162
rect 511 14 545 30
rect 607 146 641 162
rect 607 14 641 30
rect 703 146 737 162
rect 703 14 737 30
rect 799 146 833 162
rect 799 14 833 30
rect 895 146 929 162
rect 895 14 929 30
rect 991 146 1025 162
rect 991 14 1025 30
rect 1087 146 1121 162
rect 1087 14 1121 30
rect 1183 146 1217 162
rect 1183 14 1217 30
rect 1279 146 1313 162
rect 1279 14 1313 30
rect -1313 -74 -1279 -58
rect -1313 -206 -1279 -190
rect -1217 -74 -1183 -58
rect -1217 -206 -1183 -190
rect -1121 -74 -1087 -58
rect -1121 -206 -1087 -190
rect -1025 -74 -991 -58
rect -1025 -206 -991 -190
rect -929 -74 -895 -58
rect -929 -206 -895 -190
rect -833 -74 -799 -58
rect -833 -206 -799 -190
rect -737 -74 -703 -58
rect -737 -206 -703 -190
rect -641 -74 -607 -58
rect -641 -206 -607 -190
rect -545 -74 -511 -58
rect -545 -206 -511 -190
rect -449 -74 -415 -58
rect -449 -206 -415 -190
rect -353 -74 -319 -58
rect -353 -206 -319 -190
rect -257 -74 -223 -58
rect -257 -206 -223 -190
rect -161 -74 -127 -58
rect -161 -206 -127 -190
rect -65 -74 -31 -58
rect -65 -206 -31 -190
rect 31 -74 65 -58
rect 31 -206 65 -190
rect 127 -74 161 -58
rect 127 -206 161 -190
rect 223 -74 257 -58
rect 223 -206 257 -190
rect 319 -74 353 -58
rect 319 -206 353 -190
rect 415 -74 449 -58
rect 415 -206 449 -190
rect 511 -74 545 -58
rect 511 -206 545 -190
rect 607 -74 641 -58
rect 607 -206 641 -190
rect 703 -74 737 -58
rect 703 -206 737 -190
rect 799 -74 833 -58
rect 799 -206 833 -190
rect 895 -74 929 -58
rect 895 -206 929 -190
rect 991 -74 1025 -58
rect 991 -206 1025 -190
rect 1087 -74 1121 -58
rect 1087 -206 1121 -190
rect 1183 -74 1217 -58
rect 1183 -206 1217 -190
rect 1279 -74 1313 -58
rect 1279 -206 1313 -190
rect -1427 -327 -1393 -265
rect -1299 -283 -1283 -249
rect -1249 -283 -1233 -249
rect -1167 -283 -1151 -249
rect -1057 -283 -1041 -249
rect -975 -283 -959 -249
rect -289 -283 -273 -249
rect -207 -283 -191 -249
rect 1247 -283 1263 -249
rect 1393 -327 1427 -265
rect -1427 -361 -1331 -327
rect 1331 -361 1427 -327
<< viali >>
rect -1313 30 -1279 146
rect -1217 30 -1183 146
rect -1121 30 -1087 146
rect -1025 30 -991 146
rect -929 30 -895 146
rect -833 30 -799 146
rect -737 30 -703 146
rect -641 30 -607 146
rect -545 30 -511 146
rect -449 30 -415 146
rect -353 30 -319 146
rect -257 30 -223 146
rect -161 30 -127 146
rect -65 30 -31 146
rect 31 30 65 146
rect 127 30 161 146
rect 223 30 257 146
rect 319 30 353 146
rect 415 30 449 146
rect 511 30 545 146
rect 607 30 641 146
rect 703 30 737 146
rect 799 30 833 146
rect 895 30 929 146
rect 991 30 1025 146
rect 1087 30 1121 146
rect 1183 30 1217 146
rect 1279 30 1313 146
rect -1313 -190 -1279 -74
rect -1217 -190 -1183 -74
rect -1121 -190 -1087 -74
rect -1025 -190 -991 -74
rect -929 -190 -895 -74
rect -833 -190 -799 -74
rect -737 -190 -703 -74
rect -641 -190 -607 -74
rect -545 -190 -511 -74
rect -449 -190 -415 -74
rect -353 -190 -319 -74
rect -257 -190 -223 -74
rect -161 -190 -127 -74
rect -65 -190 -31 -74
rect 31 -190 65 -74
rect 127 -190 161 -74
rect 223 -190 257 -74
rect 319 -190 353 -74
rect 415 -190 449 -74
rect 511 -190 545 -74
rect 607 -190 641 -74
rect 703 -190 737 -74
rect 799 -190 833 -74
rect 895 -190 929 -74
rect 991 -190 1025 -74
rect 1087 -190 1121 -74
rect 1183 -190 1217 -74
rect 1279 -190 1313 -74
rect -1283 -283 -1249 -249
rect -1151 -283 -1057 -249
rect -959 -283 -289 -249
rect -191 -283 1247 -249
<< metal1 >>
rect -1319 146 -1273 158
rect -1319 30 -1313 146
rect -1279 30 -1273 146
rect -1319 18 -1273 30
rect -1223 146 -1177 158
rect -1223 30 -1217 146
rect -1183 30 -1177 146
rect -1223 18 -1177 30
rect -1127 146 -1081 158
rect -1127 30 -1121 146
rect -1087 30 -1081 146
rect -1127 18 -1081 30
rect -1031 146 -985 158
rect -1031 30 -1025 146
rect -991 30 -985 146
rect -1031 18 -985 30
rect -935 146 -889 158
rect -935 30 -929 146
rect -895 30 -889 146
rect -935 18 -889 30
rect -839 146 -793 158
rect -839 30 -833 146
rect -799 30 -793 146
rect -839 18 -793 30
rect -743 146 -697 158
rect -743 30 -737 146
rect -703 30 -697 146
rect -743 18 -697 30
rect -647 146 -601 158
rect -647 30 -641 146
rect -607 30 -601 146
rect -647 18 -601 30
rect -551 146 -505 158
rect -551 30 -545 146
rect -511 30 -505 146
rect -551 18 -505 30
rect -455 146 -409 158
rect -455 30 -449 146
rect -415 30 -409 146
rect -455 18 -409 30
rect -359 146 -313 158
rect -359 30 -353 146
rect -319 30 -313 146
rect -359 18 -313 30
rect -263 146 -217 158
rect -263 30 -257 146
rect -223 30 -217 146
rect -263 18 -217 30
rect -167 146 -121 158
rect -167 30 -161 146
rect -127 30 -121 146
rect -167 18 -121 30
rect -71 146 -25 158
rect -71 30 -65 146
rect -31 30 -25 146
rect -71 18 -25 30
rect 25 146 71 158
rect 25 30 31 146
rect 65 30 71 146
rect 25 18 71 30
rect 121 146 167 158
rect 121 30 127 146
rect 161 30 167 146
rect 121 18 167 30
rect 217 146 263 158
rect 217 30 223 146
rect 257 30 263 146
rect 217 18 263 30
rect 313 146 359 158
rect 313 30 319 146
rect 353 30 359 146
rect 313 18 359 30
rect 409 146 455 158
rect 409 30 415 146
rect 449 30 455 146
rect 409 18 455 30
rect 505 146 551 158
rect 505 30 511 146
rect 545 30 551 146
rect 505 18 551 30
rect 601 146 647 158
rect 601 30 607 146
rect 641 30 647 146
rect 601 18 647 30
rect 697 146 743 158
rect 697 30 703 146
rect 737 30 743 146
rect 697 18 743 30
rect 793 146 839 158
rect 793 30 799 146
rect 833 30 839 146
rect 793 18 839 30
rect 889 146 935 158
rect 889 30 895 146
rect 929 30 935 146
rect 889 18 935 30
rect 985 146 1031 158
rect 985 30 991 146
rect 1025 30 1031 146
rect 985 18 1031 30
rect 1081 146 1127 158
rect 1081 30 1087 146
rect 1121 30 1127 146
rect 1081 18 1127 30
rect 1177 146 1223 158
rect 1177 30 1183 146
rect 1217 30 1223 146
rect 1177 18 1223 30
rect 1273 146 1319 158
rect 1273 30 1279 146
rect 1313 30 1319 146
rect 1273 18 1319 30
rect -1319 -74 -1273 -62
rect -1319 -190 -1313 -74
rect -1279 -190 -1273 -74
rect -1319 -202 -1273 -190
rect -1223 -74 -1177 -62
rect -1223 -190 -1217 -74
rect -1183 -190 -1177 -74
rect -1223 -202 -1177 -190
rect -1127 -74 -1081 -62
rect -1127 -190 -1121 -74
rect -1087 -190 -1081 -74
rect -1127 -202 -1081 -190
rect -1031 -74 -985 -62
rect -1031 -190 -1025 -74
rect -991 -190 -985 -74
rect -1031 -202 -985 -190
rect -935 -74 -889 -62
rect -935 -190 -929 -74
rect -895 -190 -889 -74
rect -935 -202 -889 -190
rect -839 -74 -793 -62
rect -839 -190 -833 -74
rect -799 -190 -793 -74
rect -839 -202 -793 -190
rect -743 -74 -697 -62
rect -743 -190 -737 -74
rect -703 -190 -697 -74
rect -743 -202 -697 -190
rect -647 -74 -601 -62
rect -647 -190 -641 -74
rect -607 -190 -601 -74
rect -647 -202 -601 -190
rect -551 -74 -505 -62
rect -551 -190 -545 -74
rect -511 -190 -505 -74
rect -551 -202 -505 -190
rect -455 -74 -409 -62
rect -455 -190 -449 -74
rect -415 -190 -409 -74
rect -455 -202 -409 -190
rect -359 -74 -313 -62
rect -359 -190 -353 -74
rect -319 -190 -313 -74
rect -359 -202 -313 -190
rect -263 -74 -217 -62
rect -263 -190 -257 -74
rect -223 -190 -217 -74
rect -263 -202 -217 -190
rect -167 -74 -121 -62
rect -167 -190 -161 -74
rect -127 -190 -121 -74
rect -167 -202 -121 -190
rect -71 -74 -25 -62
rect -71 -190 -65 -74
rect -31 -190 -25 -74
rect -71 -202 -25 -190
rect 25 -74 71 -62
rect 25 -190 31 -74
rect 65 -190 71 -74
rect 25 -202 71 -190
rect 121 -74 167 -62
rect 121 -190 127 -74
rect 161 -190 167 -74
rect 121 -202 167 -190
rect 217 -74 263 -62
rect 217 -190 223 -74
rect 257 -190 263 -74
rect 217 -202 263 -190
rect 313 -74 359 -62
rect 313 -190 319 -74
rect 353 -190 359 -74
rect 313 -202 359 -190
rect 409 -74 455 -62
rect 409 -190 415 -74
rect 449 -190 455 -74
rect 409 -202 455 -190
rect 505 -74 551 -62
rect 505 -190 511 -74
rect 545 -190 551 -74
rect 505 -202 551 -190
rect 601 -74 647 -62
rect 601 -190 607 -74
rect 641 -190 647 -74
rect 601 -202 647 -190
rect 697 -74 743 -62
rect 697 -190 703 -74
rect 737 -190 743 -74
rect 697 -202 743 -190
rect 793 -74 839 -62
rect 793 -190 799 -74
rect 833 -190 839 -74
rect 793 -202 839 -190
rect 889 -74 935 -62
rect 889 -190 895 -74
rect 929 -190 935 -74
rect 889 -202 935 -190
rect 985 -74 1031 -62
rect 985 -190 991 -74
rect 1025 -190 1031 -74
rect 985 -202 1031 -190
rect 1081 -74 1127 -62
rect 1081 -190 1087 -74
rect 1121 -190 1127 -74
rect 1081 -202 1127 -190
rect 1177 -74 1223 -62
rect 1177 -190 1183 -74
rect 1217 -190 1223 -74
rect 1177 -202 1223 -190
rect 1273 -74 1319 -62
rect 1273 -190 1279 -74
rect 1313 -190 1319 -74
rect 1273 -202 1319 -190
rect -1295 -249 -1237 -243
rect -1295 -283 -1283 -249
rect -1249 -283 -1237 -249
rect -1295 -289 -1237 -283
rect -1167 -249 -1041 -243
rect -1167 -283 -1151 -249
rect -1057 -283 -1041 -249
rect -1167 -289 -1041 -283
rect -975 -249 -273 -243
rect -975 -283 -959 -249
rect -289 -283 -273 -249
rect -975 -289 -273 -283
rect -207 -249 1263 -243
rect -207 -283 -191 -249
rect 1247 -283 1263 -249
rect -207 -289 1263 -283
<< properties >>
string FIXED_BBOX -1410 -424 1410 424
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.7 l 0.15 m 2 nf 27 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
