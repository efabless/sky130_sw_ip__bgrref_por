magic
tech sky130A
magscale 1 2
timestamp 1718283729
<< nwell >>
rect -1101 -497 1101 497
<< mvpmos >>
rect -843 -200 -683 200
rect -625 -200 -465 200
rect -407 -200 -247 200
rect -189 -200 -29 200
rect 29 -200 189 200
rect 247 -200 407 200
rect 465 -200 625 200
rect 683 -200 843 200
<< mvpdiff >>
rect -901 188 -843 200
rect -901 -188 -889 188
rect -855 -188 -843 188
rect -901 -200 -843 -188
rect -683 188 -625 200
rect -683 -188 -671 188
rect -637 -188 -625 188
rect -683 -200 -625 -188
rect -465 188 -407 200
rect -465 -188 -453 188
rect -419 -188 -407 188
rect -465 -200 -407 -188
rect -247 188 -189 200
rect -247 -188 -235 188
rect -201 -188 -189 188
rect -247 -200 -189 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 189 188 247 200
rect 189 -188 201 188
rect 235 -188 247 188
rect 189 -200 247 -188
rect 407 188 465 200
rect 407 -188 419 188
rect 453 -188 465 188
rect 407 -200 465 -188
rect 625 188 683 200
rect 625 -188 637 188
rect 671 -188 683 188
rect 625 -200 683 -188
rect 843 188 901 200
rect 843 -188 855 188
rect 889 -188 901 188
rect 843 -200 901 -188
<< mvpdiffc >>
rect -889 -188 -855 188
rect -671 -188 -637 188
rect -453 -188 -419 188
rect -235 -188 -201 188
rect -17 -188 17 188
rect 201 -188 235 188
rect 419 -188 453 188
rect 637 -188 671 188
rect 855 -188 889 188
<< mvnsubdiff >>
rect -1035 419 1035 431
rect -1035 385 -927 419
rect 927 385 1035 419
rect -1035 373 1035 385
rect -1035 323 -977 373
rect -1035 -323 -1023 323
rect -989 -323 -977 323
rect 977 323 1035 373
rect -1035 -373 -977 -323
rect 977 -323 989 323
rect 1023 -323 1035 323
rect 977 -373 1035 -323
rect -1035 -385 1035 -373
rect -1035 -419 -927 -385
rect 927 -419 1035 -385
rect -1035 -431 1035 -419
<< mvnsubdiffcont >>
rect -927 385 927 419
rect -1023 -323 -989 323
rect 989 -323 1023 323
rect -927 -419 927 -385
<< poly >>
rect -843 281 -683 297
rect -843 247 -827 281
rect -699 247 -683 281
rect -843 200 -683 247
rect -625 281 -465 297
rect -625 247 -609 281
rect -481 247 -465 281
rect -625 200 -465 247
rect -407 281 -247 297
rect -407 247 -391 281
rect -263 247 -247 281
rect -407 200 -247 247
rect -189 281 -29 297
rect -189 247 -173 281
rect -45 247 -29 281
rect -189 200 -29 247
rect 29 281 189 297
rect 29 247 45 281
rect 173 247 189 281
rect 29 200 189 247
rect 247 281 407 297
rect 247 247 263 281
rect 391 247 407 281
rect 247 200 407 247
rect 465 281 625 297
rect 465 247 481 281
rect 609 247 625 281
rect 465 200 625 247
rect 683 281 843 297
rect 683 247 699 281
rect 827 247 843 281
rect 683 200 843 247
rect -843 -247 -683 -200
rect -843 -281 -827 -247
rect -699 -281 -683 -247
rect -843 -297 -683 -281
rect -625 -247 -465 -200
rect -625 -281 -609 -247
rect -481 -281 -465 -247
rect -625 -297 -465 -281
rect -407 -247 -247 -200
rect -407 -281 -391 -247
rect -263 -281 -247 -247
rect -407 -297 -247 -281
rect -189 -247 -29 -200
rect -189 -281 -173 -247
rect -45 -281 -29 -247
rect -189 -297 -29 -281
rect 29 -247 189 -200
rect 29 -281 45 -247
rect 173 -281 189 -247
rect 29 -297 189 -281
rect 247 -247 407 -200
rect 247 -281 263 -247
rect 391 -281 407 -247
rect 247 -297 407 -281
rect 465 -247 625 -200
rect 465 -281 481 -247
rect 609 -281 625 -247
rect 465 -297 625 -281
rect 683 -247 843 -200
rect 683 -281 699 -247
rect 827 -281 843 -247
rect 683 -297 843 -281
<< polycont >>
rect -827 247 -699 281
rect -609 247 -481 281
rect -391 247 -263 281
rect -173 247 -45 281
rect 45 247 173 281
rect 263 247 391 281
rect 481 247 609 281
rect 699 247 827 281
rect -827 -281 -699 -247
rect -609 -281 -481 -247
rect -391 -281 -263 -247
rect -173 -281 -45 -247
rect 45 -281 173 -247
rect 263 -281 391 -247
rect 481 -281 609 -247
rect 699 -281 827 -247
<< locali >>
rect -1023 385 -927 419
rect 927 385 1023 419
rect -1023 323 -989 385
rect 989 323 1023 385
rect -843 247 -827 281
rect -699 247 -683 281
rect -625 247 -609 281
rect -481 247 -465 281
rect -407 247 -391 281
rect -263 247 -247 281
rect -189 247 -173 281
rect -45 247 -29 281
rect 29 247 45 281
rect 173 247 189 281
rect 247 247 263 281
rect 391 247 407 281
rect 465 247 481 281
rect 609 247 625 281
rect 683 247 699 281
rect 827 247 843 281
rect -889 188 -855 204
rect -889 -204 -855 -188
rect -671 188 -637 204
rect -671 -204 -637 -188
rect -453 188 -419 204
rect -453 -204 -419 -188
rect -235 188 -201 204
rect -235 -204 -201 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 201 188 235 204
rect 201 -204 235 -188
rect 419 188 453 204
rect 419 -204 453 -188
rect 637 188 671 204
rect 637 -204 671 -188
rect 855 188 889 204
rect 855 -204 889 -188
rect -843 -281 -827 -247
rect -699 -281 -683 -247
rect -625 -281 -609 -247
rect -481 -281 -465 -247
rect -407 -281 -391 -247
rect -263 -281 -247 -247
rect -189 -281 -173 -247
rect -45 -281 -29 -247
rect 29 -281 45 -247
rect 173 -281 189 -247
rect 247 -281 263 -247
rect 391 -281 407 -247
rect 465 -281 481 -247
rect 609 -281 625 -247
rect 683 -281 699 -247
rect 827 -281 843 -247
rect -1023 -385 -989 -323
rect 989 -385 1023 -323
rect -1023 -419 -927 -385
rect 927 -419 1023 -385
<< viali >>
rect -827 247 -699 281
rect -609 247 -481 281
rect -391 247 -263 281
rect -173 247 -45 281
rect 45 247 173 281
rect 263 247 391 281
rect 481 247 609 281
rect 699 247 827 281
rect -889 -188 -855 188
rect -671 -188 -637 188
rect -453 -188 -419 188
rect -235 -188 -201 188
rect -17 -188 17 188
rect 201 -188 235 188
rect 419 -188 453 188
rect 637 -188 671 188
rect 855 -188 889 188
rect -827 -281 -699 -247
rect -609 -281 -481 -247
rect -391 -281 -263 -247
rect -173 -281 -45 -247
rect 45 -281 173 -247
rect 263 -281 391 -247
rect 481 -281 609 -247
rect 699 -281 827 -247
<< metal1 >>
rect -839 281 -687 287
rect -839 247 -827 281
rect -699 247 -687 281
rect -839 241 -687 247
rect -621 281 -469 287
rect -621 247 -609 281
rect -481 247 -469 281
rect -621 241 -469 247
rect -403 281 -251 287
rect -403 247 -391 281
rect -263 247 -251 281
rect -403 241 -251 247
rect -185 281 -33 287
rect -185 247 -173 281
rect -45 247 -33 281
rect -185 241 -33 247
rect 33 281 185 287
rect 33 247 45 281
rect 173 247 185 281
rect 33 241 185 247
rect 251 281 403 287
rect 251 247 263 281
rect 391 247 403 281
rect 251 241 403 247
rect 469 281 621 287
rect 469 247 481 281
rect 609 247 621 281
rect 469 241 621 247
rect 687 281 839 287
rect 687 247 699 281
rect 827 247 839 281
rect 687 241 839 247
rect -895 188 -849 200
rect -895 -188 -889 188
rect -855 -188 -849 188
rect -895 -200 -849 -188
rect -677 188 -631 200
rect -677 -188 -671 188
rect -637 -188 -631 188
rect -677 -200 -631 -188
rect -459 188 -413 200
rect -459 -188 -453 188
rect -419 -188 -413 188
rect -459 -200 -413 -188
rect -241 188 -195 200
rect -241 -188 -235 188
rect -201 -188 -195 188
rect -241 -200 -195 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 195 188 241 200
rect 195 -188 201 188
rect 235 -188 241 188
rect 195 -200 241 -188
rect 413 188 459 200
rect 413 -188 419 188
rect 453 -188 459 188
rect 413 -200 459 -188
rect 631 188 677 200
rect 631 -188 637 188
rect 671 -188 677 188
rect 631 -200 677 -188
rect 849 188 895 200
rect 849 -188 855 188
rect 889 -188 895 188
rect 849 -200 895 -188
rect -839 -247 -687 -241
rect -839 -281 -827 -247
rect -699 -281 -687 -247
rect -839 -287 -687 -281
rect -621 -247 -469 -241
rect -621 -281 -609 -247
rect -481 -281 -469 -247
rect -621 -287 -469 -281
rect -403 -247 -251 -241
rect -403 -281 -391 -247
rect -263 -281 -251 -247
rect -403 -287 -251 -281
rect -185 -247 -33 -241
rect -185 -281 -173 -247
rect -45 -281 -33 -247
rect -185 -287 -33 -281
rect 33 -247 185 -241
rect 33 -281 45 -247
rect 173 -281 185 -247
rect 33 -287 185 -281
rect 251 -247 403 -241
rect 251 -281 263 -247
rect 391 -281 403 -247
rect 251 -287 403 -281
rect 469 -247 621 -241
rect 469 -281 481 -247
rect 609 -281 621 -247
rect 469 -287 621 -281
rect 687 -247 839 -241
rect 687 -281 699 -247
rect 827 -281 839 -247
rect 687 -287 839 -281
<< properties >>
string FIXED_BBOX -1006 -402 1006 402
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2.0 l 0.8 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
