magic
tech sky130A
magscale 1 2
timestamp 1717363523
<< error_p >>
rect -29 281 29 287
rect -29 247 -17 281
rect -29 241 29 247
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -247 29 -241
rect -29 -281 -17 -247
rect -29 -287 29 -281
<< pwell >>
rect -226 -419 226 419
<< nmos >>
rect -30 109 30 209
rect -30 -209 30 -109
<< ndiff >>
rect -88 197 -30 209
rect -88 121 -76 197
rect -42 121 -30 197
rect -88 109 -30 121
rect 30 197 88 209
rect 30 121 42 197
rect 76 121 88 197
rect 30 109 88 121
rect -88 -121 -30 -109
rect -88 -197 -76 -121
rect -42 -197 -30 -121
rect -88 -209 -30 -197
rect 30 -121 88 -109
rect 30 -197 42 -121
rect 76 -197 88 -121
rect 30 -209 88 -197
<< ndiffc >>
rect -76 121 -42 197
rect 42 121 76 197
rect -76 -197 -42 -121
rect 42 -197 76 -121
<< psubdiff >>
rect -190 349 -94 383
rect 94 349 190 383
rect -190 287 -156 349
rect 156 287 190 349
rect -190 -349 -156 -287
rect 156 -349 190 -287
rect -190 -383 -94 -349
rect 94 -383 190 -349
<< psubdiffcont >>
rect -94 349 94 383
rect -190 -287 -156 287
rect 156 -287 190 287
rect -94 -383 94 -349
<< poly >>
rect -33 281 33 297
rect -33 247 -17 281
rect 17 247 33 281
rect -33 231 33 247
rect -30 209 30 231
rect -30 87 30 109
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -30 -109 30 -87
rect -30 -231 30 -209
rect -33 -247 33 -231
rect -33 -281 -17 -247
rect 17 -281 33 -247
rect -33 -297 33 -281
<< polycont >>
rect -17 247 17 281
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -281 17 -247
<< locali >>
rect -190 349 -94 383
rect 94 349 190 383
rect -190 287 -156 349
rect 156 287 190 349
rect -33 247 -17 281
rect 17 247 33 281
rect -76 197 -42 213
rect -76 105 -42 121
rect 42 197 76 213
rect 42 105 76 121
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -76 -121 -42 -105
rect -76 -213 -42 -197
rect 42 -121 76 -105
rect 42 -213 76 -197
rect -33 -281 -17 -247
rect 17 -281 33 -247
rect -190 -349 -156 -287
rect 156 -349 190 -287
rect -190 -383 -94 -349
rect 94 -383 190 -349
<< viali >>
rect -17 247 17 281
rect -76 121 -42 197
rect 42 121 76 197
rect -17 37 17 71
rect -17 -71 17 -37
rect -76 -197 -42 -121
rect 42 -197 76 -121
rect -17 -281 17 -247
<< metal1 >>
rect -29 281 29 287
rect -29 247 -17 281
rect 17 247 29 281
rect -29 241 29 247
rect -82 197 -36 209
rect -82 121 -76 197
rect -42 121 -36 197
rect -82 109 -36 121
rect 36 197 82 209
rect 36 121 42 197
rect 76 121 82 197
rect 36 109 82 121
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -82 -121 -36 -109
rect -82 -197 -76 -121
rect -42 -197 -36 -121
rect -82 -209 -36 -197
rect 36 -121 82 -109
rect 36 -197 42 -121
rect 76 -197 82 -121
rect 36 -209 82 -197
rect -29 -247 29 -241
rect -29 -281 -17 -247
rect 17 -281 29 -247
rect -29 -287 29 -281
<< properties >>
string FIXED_BBOX -173 -366 173 366
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.3 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
