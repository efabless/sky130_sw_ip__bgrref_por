magic
tech sky130A
timestamp 1717363523
<< pwell >>
rect -139 -309 139 309
<< mvnmos >>
rect -25 -180 25 180
<< mvndiff >>
rect -54 174 -25 180
rect -54 -174 -48 174
rect -31 -174 -25 174
rect -54 -180 -25 -174
rect 25 174 54 180
rect 25 -174 31 174
rect 48 -174 54 174
rect 25 -180 54 -174
<< mvndiffc >>
rect -48 -174 -31 174
rect 31 -174 48 174
<< mvpsubdiff >>
rect -121 285 121 291
rect -121 268 -67 285
rect 67 268 121 285
rect -121 262 121 268
rect -121 237 -92 262
rect -121 -237 -115 237
rect -98 -237 -92 237
rect 92 237 121 262
rect -121 -262 -92 -237
rect 92 -237 98 237
rect 115 -237 121 237
rect 92 -262 121 -237
rect -121 -268 121 -262
rect -121 -285 -67 -268
rect 67 -285 121 -268
rect -121 -291 121 -285
<< mvpsubdiffcont >>
rect -67 268 67 285
rect -115 -237 -98 237
rect 98 -237 115 237
rect -67 -285 67 -268
<< poly >>
rect -25 216 25 224
rect -25 199 -17 216
rect 17 199 25 216
rect -25 180 25 199
rect -25 -199 25 -180
rect -25 -216 -17 -199
rect 17 -216 25 -199
rect -25 -224 25 -216
<< polycont >>
rect -17 199 17 216
rect -17 -216 17 -199
<< locali >>
rect -115 268 -67 285
rect 67 268 115 285
rect -115 237 -98 268
rect 98 237 115 268
rect -25 199 -17 216
rect 17 199 25 216
rect -48 174 -31 182
rect -48 -182 -31 -174
rect 31 174 48 182
rect 31 -182 48 -174
rect -25 -216 -17 -199
rect 17 -216 25 -199
rect -115 -268 -98 -237
rect 98 -268 115 -237
rect -115 -285 -67 -268
rect 67 -285 115 -268
<< viali >>
rect -17 199 17 216
rect -48 -174 -31 174
rect 31 -174 48 174
rect -17 -216 17 -199
<< metal1 >>
rect -23 216 23 219
rect -23 199 -17 216
rect 17 199 23 216
rect -23 196 23 199
rect -51 174 -28 180
rect -51 -174 -48 174
rect -31 -174 -28 174
rect -51 -180 -28 -174
rect 28 174 51 180
rect 28 -174 31 174
rect 48 -174 51 174
rect 28 -180 51 -174
rect -23 -199 23 -196
rect -23 -216 -17 -199
rect 17 -216 23 -199
rect -23 -219 23 -216
<< properties >>
string FIXED_BBOX -106 -276 106 276
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 3.6 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
