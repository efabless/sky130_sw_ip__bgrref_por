magic
tech sky130A
magscale 1 2
timestamp 1721073345
<< locali >>
rect 42106 -285972 42347 -285968
rect 42106 -286006 42121 -285972
rect 42329 -286006 42347 -285972
rect 42106 -286013 42347 -286006
rect 42386 -285999 42442 -285986
rect 41522 -286065 41756 -286053
rect 41522 -286116 41537 -286065
rect 41740 -286116 41756 -286065
rect 41522 -286129 41756 -286116
rect 41870 -286068 42167 -286060
rect 41870 -286114 41890 -286068
rect 42143 -286114 42167 -286068
rect 41870 -286121 42167 -286114
rect 42386 -286202 42394 -285999
rect 42430 -286202 42442 -285999
rect 42545 -286028 42597 -286025
rect 42545 -286062 42554 -286028
rect 42588 -286062 42597 -286028
rect 42545 -286153 42597 -286062
rect 42660 -286027 42722 -286020
rect 42660 -286068 42678 -286027
rect 42713 -286068 42722 -286027
rect 42660 -286074 42722 -286068
rect 42386 -286217 42442 -286202
rect 42182 -286555 42246 -286542
rect 42182 -286744 42192 -286555
rect 42235 -286744 42246 -286555
rect 42182 -286753 42246 -286744
rect 42398 -286704 42464 -286691
rect 41250 -286780 41496 -286768
rect 41250 -286829 41265 -286780
rect 41481 -286829 41496 -286780
rect 41250 -286842 41496 -286829
rect 42398 -286888 42410 -286704
rect 42453 -286888 42464 -286704
rect 42398 -286903 42464 -286888
rect 42574 -286764 42626 -286690
rect 42574 -286890 42577 -286764
rect 42623 -286890 42626 -286764
rect 42777 -286768 42824 -286761
rect 42777 -286848 42780 -286768
rect 42821 -286848 42824 -286768
rect 42777 -286854 42824 -286848
rect 42574 -286899 42626 -286890
<< viali >>
rect 42121 -286006 42329 -285972
rect 41537 -286116 41740 -286065
rect 41890 -286114 42143 -286068
rect 42394 -286202 42430 -285999
rect 42554 -286062 42588 -286028
rect 42678 -286068 42713 -286027
rect 44505 -286342 44556 -286190
rect 42192 -286744 42235 -286555
rect 41265 -286829 41481 -286780
rect 42410 -286888 42453 -286704
rect 44325 -286704 44376 -286552
rect 42577 -286890 42623 -286764
rect 42780 -286848 42821 -286768
<< metal1 >>
rect 40255 -285844 44687 -285733
rect 40846 -286395 40963 -285897
rect 41015 -285931 44687 -285844
rect 42106 -285967 42347 -285966
rect 41363 -285972 42347 -285967
rect 41363 -286004 42121 -285972
rect 42106 -286006 42121 -286004
rect 42329 -286006 42347 -285972
rect 42106 -286013 42347 -286006
rect 42383 -285999 42442 -285986
rect 41522 -286065 41756 -286053
rect 41522 -286116 41537 -286065
rect 41740 -286116 41756 -286065
rect 41522 -286129 41756 -286116
rect 41870 -286068 42167 -286060
rect 41870 -286114 41890 -286068
rect 42143 -286114 42167 -286068
rect 41870 -286121 42167 -286114
rect 42383 -286202 42394 -285999
rect 42430 -286202 42442 -285999
rect 42538 -286028 42605 -286019
rect 42538 -286062 42554 -286028
rect 42588 -286062 42605 -286028
rect 42538 -286162 42605 -286062
rect 42661 -286027 42728 -286015
rect 42661 -286068 42678 -286027
rect 42713 -286068 42728 -286027
rect 42661 -286074 42728 -286068
rect 42383 -286217 42442 -286202
rect 44493 -286190 44569 -286179
rect 44493 -286342 44505 -286190
rect 44556 -286236 44569 -286190
rect 44556 -286276 44741 -286236
rect 44556 -286342 44569 -286276
rect 44493 -286356 44569 -286342
rect 40846 -286512 44741 -286395
rect 42182 -286555 42246 -286542
rect 40960 -286670 41089 -286632
rect 41051 -286865 41089 -286670
rect 42182 -286744 42192 -286555
rect 42235 -286744 42246 -286555
rect 44313 -286552 44389 -286541
rect 42388 -286704 42464 -286691
rect 42388 -286711 42410 -286704
rect 42182 -286758 42246 -286744
rect 41250 -286780 41496 -286768
rect 41250 -286829 41265 -286780
rect 41481 -286829 41496 -286780
rect 41250 -286836 41496 -286829
rect 42398 -286865 42410 -286711
rect 41051 -286888 42410 -286865
rect 42453 -286888 42464 -286704
rect 41051 -286903 42464 -286888
rect 42566 -286764 42633 -286683
rect 44313 -286704 44325 -286552
rect 44376 -286596 44389 -286552
rect 44376 -286636 44741 -286596
rect 44376 -286704 44389 -286636
rect 44313 -286718 44389 -286704
rect 42566 -286890 42577 -286764
rect 42623 -286890 42633 -286764
rect 42768 -286768 42833 -286751
rect 42768 -286848 42780 -286768
rect 42821 -286848 42833 -286768
rect 42768 -286863 42833 -286848
rect 42566 -286907 42633 -286890
rect 40248 -287162 44680 -286945
<< metal2 >>
rect 42193 -285969 42701 -285934
rect 40878 -286642 40952 -286567
rect 41363 -286788 41400 -286004
rect 41614 -287190 41656 -286105
rect 41974 -287179 42016 -286094
rect 42193 -286656 42228 -285969
rect 42666 -286055 42701 -285969
rect 42382 -286819 42437 -286087
rect 42560 -286394 42601 -286084
rect 42560 -286427 42824 -286394
rect 42560 -286435 42826 -286427
rect 42579 -287173 42620 -286873
rect 42785 -287172 42826 -286435
use por_via_2cut  por_via_2cut_185
timestamp 1718283729
transform 0 1 50703 -1 0 -270664
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_188
timestamp 1718283729
transform 1 0 24776 0 1 -278754
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_191
timestamp 1718283729
transform 0 1 50310 -1 0 -269996
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_192
timestamp 1718283729
transform 0 1 50314 -1 0 -270597
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_193
timestamp 1718283729
transform 0 1 50113 -1 0 -270483
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_194
timestamp 1718283729
transform -1 0 57529 0 -1 -294702
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_195
timestamp 1718283729
transform 0 1 50472 -1 0 -269926
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_196
timestamp 1718283729
transform -1 0 58876 0 -1 -293941
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_197
timestamp 1718283729
transform -1 0 57582 0 -1 -293900
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_198
timestamp 1718283729
transform -1 0 57799 0 -1 -293991
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_199
timestamp 1718283729
transform -1 0 58166 0 -1 -293991
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_201
timestamp 1718283729
transform 0 1 50500 -1 0 -270670
box 16088 -7932 16222 -7868
use sky130_fd_sc_ls__buf_8  sky130_fd_sc_ls__buf_8_0 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1715205430
transform 1 0 41217 0 1 -287116
box -38 -49 1190 715
use sky130_fd_sc_ls__decap_4  sky130_fd_sc_ls__decap_4_0 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1715205430
transform 1 0 41121 0 -1 -285784
box -38 -49 422 715
use sky130_fd_sc_ls__dfrtn_1  sky130_fd_sc_ls__dfrtn_1_0 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1715205430
transform 1 0 42369 0 -1 -285784
box -38 -49 2246 715
use sky130_fd_sc_ls__dfrtp_1  sky130_fd_sc_ls__dfrtp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1715205430
transform 1 0 42369 0 1 -287116
box -38 -49 2246 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  sky130_fd_sc_ls__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1715205430
transform 1 0 41505 0 -1 -285784
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  sky130_fd_sc_ls__tapvpwrvgnd_1_1
timestamp 1715205430
transform 1 0 44577 0 -1 -285784
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  sky130_fd_sc_ls__tapvpwrvgnd_1_2
timestamp 1715205430
transform 1 0 41121 0 1 -287116
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  sky130_fd_sc_ls__tapvpwrvgnd_1_3
timestamp 1715205430
transform 1 0 44577 0 1 -287116
box -38 -49 134 715
use sky130_fd_sc_ls__xor2_1  sky130_fd_sc_ls__xor2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1715205430
transform 1 0 41601 0 -1 -285784
box -38 -49 806 715
use TieH_1p8  TieH_1p8_0
timestamp 1718283729
transform 1 0 39912 0 1 -286191
box 346 -837 1050 296
<< end >>
