magic
tech sky130A
magscale 1 2
timestamp 1717363523
<< pwell >>
rect -296 -1955 296 1955
<< nmos >>
rect -100 1345 100 1745
rect -100 727 100 1127
rect -100 109 100 509
rect -100 -509 100 -109
rect -100 -1127 100 -727
rect -100 -1745 100 -1345
<< ndiff >>
rect -158 1733 -100 1745
rect -158 1357 -146 1733
rect -112 1357 -100 1733
rect -158 1345 -100 1357
rect 100 1733 158 1745
rect 100 1357 112 1733
rect 146 1357 158 1733
rect 100 1345 158 1357
rect -158 1115 -100 1127
rect -158 739 -146 1115
rect -112 739 -100 1115
rect -158 727 -100 739
rect 100 1115 158 1127
rect 100 739 112 1115
rect 146 739 158 1115
rect 100 727 158 739
rect -158 497 -100 509
rect -158 121 -146 497
rect -112 121 -100 497
rect -158 109 -100 121
rect 100 497 158 509
rect 100 121 112 497
rect 146 121 158 497
rect 100 109 158 121
rect -158 -121 -100 -109
rect -158 -497 -146 -121
rect -112 -497 -100 -121
rect -158 -509 -100 -497
rect 100 -121 158 -109
rect 100 -497 112 -121
rect 146 -497 158 -121
rect 100 -509 158 -497
rect -158 -739 -100 -727
rect -158 -1115 -146 -739
rect -112 -1115 -100 -739
rect -158 -1127 -100 -1115
rect 100 -739 158 -727
rect 100 -1115 112 -739
rect 146 -1115 158 -739
rect 100 -1127 158 -1115
rect -158 -1357 -100 -1345
rect -158 -1733 -146 -1357
rect -112 -1733 -100 -1357
rect -158 -1745 -100 -1733
rect 100 -1357 158 -1345
rect 100 -1733 112 -1357
rect 146 -1733 158 -1357
rect 100 -1745 158 -1733
<< ndiffc >>
rect -146 1357 -112 1733
rect 112 1357 146 1733
rect -146 739 -112 1115
rect 112 739 146 1115
rect -146 121 -112 497
rect 112 121 146 497
rect -146 -497 -112 -121
rect 112 -497 146 -121
rect -146 -1115 -112 -739
rect 112 -1115 146 -739
rect -146 -1733 -112 -1357
rect 112 -1733 146 -1357
<< psubdiff >>
rect -260 1885 -164 1919
rect 164 1885 260 1919
rect -260 1823 -226 1885
rect 226 1823 260 1885
rect -260 -1885 -226 -1823
rect 226 -1885 260 -1823
rect -260 -1919 -164 -1885
rect 164 -1919 260 -1885
<< psubdiffcont >>
rect -164 1885 164 1919
rect -260 -1823 -226 1823
rect 226 -1823 260 1823
rect -164 -1919 164 -1885
<< poly >>
rect -100 1817 100 1833
rect -100 1783 -84 1817
rect 84 1783 100 1817
rect -100 1745 100 1783
rect -100 1307 100 1345
rect -100 1273 -84 1307
rect 84 1273 100 1307
rect -100 1257 100 1273
rect -100 1199 100 1215
rect -100 1165 -84 1199
rect 84 1165 100 1199
rect -100 1127 100 1165
rect -100 689 100 727
rect -100 655 -84 689
rect 84 655 100 689
rect -100 639 100 655
rect -100 581 100 597
rect -100 547 -84 581
rect 84 547 100 581
rect -100 509 100 547
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -109 100 -71
rect -100 -547 100 -509
rect -100 -581 -84 -547
rect 84 -581 100 -547
rect -100 -597 100 -581
rect -100 -655 100 -639
rect -100 -689 -84 -655
rect 84 -689 100 -655
rect -100 -727 100 -689
rect -100 -1165 100 -1127
rect -100 -1199 -84 -1165
rect 84 -1199 100 -1165
rect -100 -1215 100 -1199
rect -100 -1273 100 -1257
rect -100 -1307 -84 -1273
rect 84 -1307 100 -1273
rect -100 -1345 100 -1307
rect -100 -1783 100 -1745
rect -100 -1817 -84 -1783
rect 84 -1817 100 -1783
rect -100 -1833 100 -1817
<< polycont >>
rect -84 1783 84 1817
rect -84 1273 84 1307
rect -84 1165 84 1199
rect -84 655 84 689
rect -84 547 84 581
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -581 84 -547
rect -84 -689 84 -655
rect -84 -1199 84 -1165
rect -84 -1307 84 -1273
rect -84 -1817 84 -1783
<< locali >>
rect -260 1885 -164 1919
rect 164 1885 260 1919
rect -260 1823 -226 1885
rect 226 1823 260 1885
rect -100 1783 -84 1817
rect 84 1783 100 1817
rect -146 1733 -112 1749
rect -146 1341 -112 1357
rect 112 1733 146 1749
rect 112 1341 146 1357
rect -100 1273 -84 1307
rect 84 1273 100 1307
rect -100 1165 -84 1199
rect 84 1165 100 1199
rect -146 1115 -112 1131
rect -146 723 -112 739
rect 112 1115 146 1131
rect 112 723 146 739
rect -100 655 -84 689
rect 84 655 100 689
rect -100 547 -84 581
rect 84 547 100 581
rect -146 497 -112 513
rect -146 105 -112 121
rect 112 497 146 513
rect 112 105 146 121
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -121 -112 -105
rect -146 -513 -112 -497
rect 112 -121 146 -105
rect 112 -513 146 -497
rect -100 -581 -84 -547
rect 84 -581 100 -547
rect -100 -689 -84 -655
rect 84 -689 100 -655
rect -146 -739 -112 -723
rect -146 -1131 -112 -1115
rect 112 -739 146 -723
rect 112 -1131 146 -1115
rect -100 -1199 -84 -1165
rect 84 -1199 100 -1165
rect -100 -1307 -84 -1273
rect 84 -1307 100 -1273
rect -146 -1357 -112 -1341
rect -146 -1749 -112 -1733
rect 112 -1357 146 -1341
rect 112 -1749 146 -1733
rect -100 -1817 -84 -1783
rect 84 -1817 100 -1783
rect -260 -1885 -226 -1823
rect 226 -1885 260 -1823
rect -260 -1919 -164 -1885
rect 164 -1919 260 -1885
<< viali >>
rect -84 1783 84 1817
rect -146 1357 -112 1733
rect 112 1357 146 1733
rect -84 1273 84 1307
rect -84 1165 84 1199
rect -146 739 -112 1115
rect 112 739 146 1115
rect -84 655 84 689
rect -84 547 84 581
rect -146 121 -112 497
rect 112 121 146 497
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -497 -112 -121
rect 112 -497 146 -121
rect -84 -581 84 -547
rect -84 -689 84 -655
rect -146 -1115 -112 -739
rect 112 -1115 146 -739
rect -84 -1199 84 -1165
rect -84 -1307 84 -1273
rect -146 -1733 -112 -1357
rect 112 -1733 146 -1357
rect -84 -1817 84 -1783
<< metal1 >>
rect -96 1817 96 1823
rect -96 1783 -84 1817
rect 84 1783 96 1817
rect -96 1777 96 1783
rect -152 1733 -106 1745
rect -152 1357 -146 1733
rect -112 1357 -106 1733
rect -152 1345 -106 1357
rect 106 1733 152 1745
rect 106 1357 112 1733
rect 146 1357 152 1733
rect 106 1345 152 1357
rect -96 1307 96 1313
rect -96 1273 -84 1307
rect 84 1273 96 1307
rect -96 1267 96 1273
rect -96 1199 96 1205
rect -96 1165 -84 1199
rect 84 1165 96 1199
rect -96 1159 96 1165
rect -152 1115 -106 1127
rect -152 739 -146 1115
rect -112 739 -106 1115
rect -152 727 -106 739
rect 106 1115 152 1127
rect 106 739 112 1115
rect 146 739 152 1115
rect 106 727 152 739
rect -96 689 96 695
rect -96 655 -84 689
rect 84 655 96 689
rect -96 649 96 655
rect -96 581 96 587
rect -96 547 -84 581
rect 84 547 96 581
rect -96 541 96 547
rect -152 497 -106 509
rect -152 121 -146 497
rect -112 121 -106 497
rect -152 109 -106 121
rect 106 497 152 509
rect 106 121 112 497
rect 146 121 152 497
rect 106 109 152 121
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -121 -106 -109
rect -152 -497 -146 -121
rect -112 -497 -106 -121
rect -152 -509 -106 -497
rect 106 -121 152 -109
rect 106 -497 112 -121
rect 146 -497 152 -121
rect 106 -509 152 -497
rect -96 -547 96 -541
rect -96 -581 -84 -547
rect 84 -581 96 -547
rect -96 -587 96 -581
rect -96 -655 96 -649
rect -96 -689 -84 -655
rect 84 -689 96 -655
rect -96 -695 96 -689
rect -152 -739 -106 -727
rect -152 -1115 -146 -739
rect -112 -1115 -106 -739
rect -152 -1127 -106 -1115
rect 106 -739 152 -727
rect 106 -1115 112 -739
rect 146 -1115 152 -739
rect 106 -1127 152 -1115
rect -96 -1165 96 -1159
rect -96 -1199 -84 -1165
rect 84 -1199 96 -1165
rect -96 -1205 96 -1199
rect -96 -1273 96 -1267
rect -96 -1307 -84 -1273
rect 84 -1307 96 -1273
rect -96 -1313 96 -1307
rect -152 -1357 -106 -1345
rect -152 -1733 -146 -1357
rect -112 -1733 -106 -1357
rect -152 -1745 -106 -1733
rect 106 -1357 152 -1345
rect 106 -1733 112 -1357
rect 146 -1733 152 -1357
rect 106 -1745 152 -1733
rect -96 -1783 96 -1777
rect -96 -1817 -84 -1783
rect 84 -1817 96 -1783
rect -96 -1823 96 -1817
<< properties >>
string FIXED_BBOX -243 -1902 243 1902
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.0 l 1.0 m 6 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
