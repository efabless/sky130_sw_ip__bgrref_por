magic
tech sky130A
magscale 1 2
timestamp 1717363523
<< metal4 >>
rect -1949 5239 1949 5280
rect -1949 1961 1693 5239
rect 1929 1961 1949 5239
rect -1949 1920 1949 1961
rect -1949 1639 1949 1680
rect -1949 -1639 1693 1639
rect 1929 -1639 1949 1639
rect -1949 -1680 1949 -1639
rect -1949 -1961 1949 -1920
rect -1949 -5239 1693 -1961
rect 1929 -5239 1949 -1961
rect -1949 -5280 1949 -5239
<< via4 >>
rect 1693 1961 1929 5239
rect 1693 -1639 1929 1639
rect 1693 -5239 1929 -1961
<< mimcap2 >>
rect -1869 5160 1331 5200
rect -1869 2040 -1829 5160
rect 1291 2040 1331 5160
rect -1869 2000 1331 2040
rect -1869 1560 1331 1600
rect -1869 -1560 -1829 1560
rect 1291 -1560 1331 1560
rect -1869 -1600 1331 -1560
rect -1869 -2040 1331 -2000
rect -1869 -5160 -1829 -2040
rect 1291 -5160 1331 -2040
rect -1869 -5200 1331 -5160
<< mimcap2contact >>
rect -1829 2040 1291 5160
rect -1829 -1560 1291 1560
rect -1829 -5160 1291 -2040
<< metal5 >>
rect -429 5184 -109 5400
rect 1651 5239 1971 5400
rect -1853 5160 1315 5184
rect -1853 2040 -1829 5160
rect 1291 2040 1315 5160
rect -1853 2016 1315 2040
rect -429 1584 -109 2016
rect 1651 1961 1693 5239
rect 1929 1961 1971 5239
rect 1651 1639 1971 1961
rect -1853 1560 1315 1584
rect -1853 -1560 -1829 1560
rect 1291 -1560 1315 1560
rect -1853 -1584 1315 -1560
rect -429 -2016 -109 -1584
rect 1651 -1639 1693 1639
rect 1929 -1639 1971 1639
rect 1651 -1961 1971 -1639
rect -1853 -2040 1315 -2016
rect -1853 -5160 -1829 -2040
rect 1291 -5160 1315 -2040
rect -1853 -5184 1315 -5160
rect -429 -5400 -109 -5184
rect 1651 -5239 1693 -1961
rect 1929 -5239 1971 -1961
rect 1651 -5400 1971 -5239
<< properties >>
string FIXED_BBOX -1949 1920 1411 5280
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 16.0 l 16.0 val 524.159 carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
