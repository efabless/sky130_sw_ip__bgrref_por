magic
tech sky130A
magscale 1 2
timestamp 1717438235
<< metal3 >>
rect -9362 9272 -5890 9300
rect -9362 6248 -5974 9272
rect -5910 6248 -5890 9272
rect -9362 6220 -5890 6248
rect -5064 9272 -1592 9300
rect -5064 6248 -1676 9272
rect -1612 6248 -1592 9272
rect -5064 6220 -1592 6248
rect -766 9272 2706 9300
rect -766 6248 2622 9272
rect 2686 6248 2706 9272
rect -766 6220 2706 6248
rect 3532 9272 7004 9300
rect 3532 6248 6920 9272
rect 6984 6248 7004 9272
rect 3532 6220 7004 6248
rect -9362 5672 -5890 5700
rect -9362 2648 -5974 5672
rect -5910 2648 -5890 5672
rect -9362 2620 -5890 2648
rect -5064 5672 -1592 5700
rect -5064 2648 -1676 5672
rect -1612 2648 -1592 5672
rect -5064 2620 -1592 2648
rect -766 5672 2706 5700
rect -766 2648 2622 5672
rect 2686 2648 2706 5672
rect -766 2620 2706 2648
rect 3532 5672 7004 5700
rect 3532 2648 6920 5672
rect 6984 2648 7004 5672
rect 3532 2620 7004 2648
rect -9362 2072 -5890 2100
rect -9362 -952 -5974 2072
rect -5910 -952 -5890 2072
rect -9362 -980 -5890 -952
rect -5064 2072 -1592 2100
rect -5064 -952 -1676 2072
rect -1612 -952 -1592 2072
rect -5064 -980 -1592 -952
rect -766 2072 2706 2100
rect -766 -952 2622 2072
rect 2686 -952 2706 2072
rect -766 -980 2706 -952
rect 3532 2072 7004 2100
rect 3532 -952 6920 2072
rect 6984 -952 7004 2072
rect 3532 -980 7004 -952
rect -9362 -1528 -5890 -1500
rect -9362 -4552 -5974 -1528
rect -5910 -4552 -5890 -1528
rect -9362 -4580 -5890 -4552
rect -5064 -1528 -1592 -1500
rect -5064 -4552 -1676 -1528
rect -1612 -4552 -1592 -1528
rect -5064 -4580 -1592 -4552
rect -766 -1528 2706 -1500
rect -766 -4552 2622 -1528
rect 2686 -4552 2706 -1528
rect -766 -4580 2706 -4552
rect 3532 -1528 7004 -1500
rect 3532 -4552 6920 -1528
rect 6984 -4552 7004 -1528
rect 3532 -4580 7004 -4552
rect -9362 -5128 -5890 -5100
rect -9362 -8152 -5974 -5128
rect -5910 -8152 -5890 -5128
rect -9362 -8180 -5890 -8152
rect -5064 -5128 -1592 -5100
rect -5064 -8152 -1676 -5128
rect -1612 -8152 -1592 -5128
rect -5064 -8180 -1592 -8152
rect -766 -5128 2706 -5100
rect -766 -8152 2622 -5128
rect 2686 -8152 2706 -5128
rect -766 -8180 2706 -8152
rect 3532 -5128 7004 -5100
rect 3532 -8152 6920 -5128
rect 6984 -8152 7004 -5128
rect 3532 -8180 7004 -8152
<< via3 >>
rect -5974 6248 -5910 9272
rect -1676 6248 -1612 9272
rect 2622 6248 2686 9272
rect 6920 6248 6984 9272
rect -5974 2648 -5910 5672
rect -1676 2648 -1612 5672
rect 2622 2648 2686 5672
rect 6920 2648 6984 5672
rect -5974 -952 -5910 2072
rect -1676 -952 -1612 2072
rect 2622 -952 2686 2072
rect 6920 -952 6984 2072
rect -5974 -4552 -5910 -1528
rect -1676 -4552 -1612 -1528
rect 2622 -4552 2686 -1528
rect 6920 -4552 6984 -1528
rect -5974 -8152 -5910 -5128
rect -1676 -8152 -1612 -5128
rect 2622 -8152 2686 -5128
rect 6920 -8152 6984 -5128
<< mimcap >>
rect -9322 9220 -6322 9260
rect -9322 6300 -9282 9220
rect -6362 6300 -6322 9220
rect -9322 6260 -6322 6300
rect -5024 9220 -2024 9260
rect -5024 6300 -4984 9220
rect -2064 6300 -2024 9220
rect -5024 6260 -2024 6300
rect -726 9220 2274 9260
rect -726 6300 -686 9220
rect 2234 6300 2274 9220
rect -726 6260 2274 6300
rect 3572 9220 6572 9260
rect 3572 6300 3612 9220
rect 6532 6300 6572 9220
rect 3572 6260 6572 6300
rect -9322 5620 -6322 5660
rect -9322 2700 -9282 5620
rect -6362 2700 -6322 5620
rect -9322 2660 -6322 2700
rect -5024 5620 -2024 5660
rect -5024 2700 -4984 5620
rect -2064 2700 -2024 5620
rect -5024 2660 -2024 2700
rect -726 5620 2274 5660
rect -726 2700 -686 5620
rect 2234 2700 2274 5620
rect -726 2660 2274 2700
rect 3572 5620 6572 5660
rect 3572 2700 3612 5620
rect 6532 2700 6572 5620
rect 3572 2660 6572 2700
rect -9322 2020 -6322 2060
rect -9322 -900 -9282 2020
rect -6362 -900 -6322 2020
rect -9322 -940 -6322 -900
rect -5024 2020 -2024 2060
rect -5024 -900 -4984 2020
rect -2064 -900 -2024 2020
rect -5024 -940 -2024 -900
rect -726 2020 2274 2060
rect -726 -900 -686 2020
rect 2234 -900 2274 2020
rect -726 -940 2274 -900
rect 3572 2020 6572 2060
rect 3572 -900 3612 2020
rect 6532 -900 6572 2020
rect 3572 -940 6572 -900
rect -9322 -1580 -6322 -1540
rect -9322 -4500 -9282 -1580
rect -6362 -4500 -6322 -1580
rect -9322 -4540 -6322 -4500
rect -5024 -1580 -2024 -1540
rect -5024 -4500 -4984 -1580
rect -2064 -4500 -2024 -1580
rect -5024 -4540 -2024 -4500
rect -726 -1580 2274 -1540
rect -726 -4500 -686 -1580
rect 2234 -4500 2274 -1580
rect -726 -4540 2274 -4500
rect 3572 -1580 6572 -1540
rect 3572 -4500 3612 -1580
rect 6532 -4500 6572 -1580
rect 3572 -4540 6572 -4500
rect -9322 -5180 -6322 -5140
rect -9322 -8100 -9282 -5180
rect -6362 -8100 -6322 -5180
rect -9322 -8140 -6322 -8100
rect -5024 -5180 -2024 -5140
rect -5024 -8100 -4984 -5180
rect -2064 -8100 -2024 -5180
rect -5024 -8140 -2024 -8100
rect -726 -5180 2274 -5140
rect -726 -8100 -686 -5180
rect 2234 -8100 2274 -5180
rect -726 -8140 2274 -8100
rect 3572 -5180 6572 -5140
rect 3572 -8100 3612 -5180
rect 6532 -8100 6572 -5180
rect 3572 -8140 6572 -8100
<< mimcapcontact >>
rect -9282 6300 -6362 9220
rect -4984 6300 -2064 9220
rect -686 6300 2234 9220
rect 3612 6300 6532 9220
rect -9282 2700 -6362 5620
rect -4984 2700 -2064 5620
rect -686 2700 2234 5620
rect 3612 2700 6532 5620
rect -9282 -900 -6362 2020
rect -4984 -900 -2064 2020
rect -686 -900 2234 2020
rect 3612 -900 6532 2020
rect -9282 -4500 -6362 -1580
rect -4984 -4500 -2064 -1580
rect -686 -4500 2234 -1580
rect 3612 -4500 6532 -1580
rect -9282 -8100 -6362 -5180
rect -4984 -8100 -2064 -5180
rect -686 -8100 2234 -5180
rect 3612 -8100 6532 -5180
<< metal4 >>
rect -7874 9221 -7770 9420
rect -5994 9272 -5890 9420
rect -9283 9220 -6361 9221
rect -9283 6300 -9282 9220
rect -6362 6300 -6361 9220
rect -9283 6299 -6361 6300
rect -7874 5621 -7770 6299
rect -5994 6248 -5974 9272
rect -5910 6248 -5890 9272
rect -3576 9221 -3472 9420
rect -1696 9272 -1592 9420
rect -4985 9220 -2063 9221
rect -4985 6300 -4984 9220
rect -2064 6300 -2063 9220
rect -4985 6299 -2063 6300
rect -5994 5672 -5890 6248
rect -9283 5620 -6361 5621
rect -9283 2700 -9282 5620
rect -6362 2700 -6361 5620
rect -9283 2699 -6361 2700
rect -7874 2021 -7770 2699
rect -5994 2648 -5974 5672
rect -5910 2648 -5890 5672
rect -3576 5621 -3472 6299
rect -1696 6248 -1676 9272
rect -1612 6248 -1592 9272
rect 722 9221 826 9420
rect 2602 9272 2706 9420
rect -687 9220 2235 9221
rect -687 6300 -686 9220
rect 2234 6300 2235 9220
rect -687 6299 2235 6300
rect -1696 5672 -1592 6248
rect -4985 5620 -2063 5621
rect -4985 2700 -4984 5620
rect -2064 2700 -2063 5620
rect -4985 2699 -2063 2700
rect -5994 2072 -5890 2648
rect -9283 2020 -6361 2021
rect -9283 -900 -9282 2020
rect -6362 -900 -6361 2020
rect -9283 -901 -6361 -900
rect -7874 -1579 -7770 -901
rect -5994 -952 -5974 2072
rect -5910 -952 -5890 2072
rect -3576 2021 -3472 2699
rect -1696 2648 -1676 5672
rect -1612 2648 -1592 5672
rect 722 5621 826 6299
rect 2602 6248 2622 9272
rect 2686 6248 2706 9272
rect 5020 9221 5124 9420
rect 6900 9272 7004 9420
rect 3611 9220 6533 9221
rect 3611 6300 3612 9220
rect 6532 6300 6533 9220
rect 3611 6299 6533 6300
rect 2602 5672 2706 6248
rect -687 5620 2235 5621
rect -687 2700 -686 5620
rect 2234 2700 2235 5620
rect -687 2699 2235 2700
rect -1696 2072 -1592 2648
rect -4985 2020 -2063 2021
rect -4985 -900 -4984 2020
rect -2064 -900 -2063 2020
rect -4985 -901 -2063 -900
rect -5994 -1528 -5890 -952
rect -9283 -1580 -6361 -1579
rect -9283 -4500 -9282 -1580
rect -6362 -4500 -6361 -1580
rect -9283 -4501 -6361 -4500
rect -7874 -5179 -7770 -4501
rect -5994 -4552 -5974 -1528
rect -5910 -4552 -5890 -1528
rect -3576 -1579 -3472 -901
rect -1696 -952 -1676 2072
rect -1612 -952 -1592 2072
rect 722 2021 826 2699
rect 2602 2648 2622 5672
rect 2686 2648 2706 5672
rect 5020 5621 5124 6299
rect 6900 6248 6920 9272
rect 6984 6248 7004 9272
rect 6900 5672 7004 6248
rect 3611 5620 6533 5621
rect 3611 2700 3612 5620
rect 6532 2700 6533 5620
rect 3611 2699 6533 2700
rect 2602 2072 2706 2648
rect -687 2020 2235 2021
rect -687 -900 -686 2020
rect 2234 -900 2235 2020
rect -687 -901 2235 -900
rect -1696 -1528 -1592 -952
rect -4985 -1580 -2063 -1579
rect -4985 -4500 -4984 -1580
rect -2064 -4500 -2063 -1580
rect -4985 -4501 -2063 -4500
rect -5994 -5128 -5890 -4552
rect -9283 -5180 -6361 -5179
rect -9283 -8100 -9282 -5180
rect -6362 -8100 -6361 -5180
rect -9283 -8101 -6361 -8100
rect -7874 -8300 -7770 -8101
rect -5994 -8152 -5974 -5128
rect -5910 -8152 -5890 -5128
rect -3576 -5179 -3472 -4501
rect -1696 -4552 -1676 -1528
rect -1612 -4552 -1592 -1528
rect 722 -1579 826 -901
rect 2602 -952 2622 2072
rect 2686 -952 2706 2072
rect 5020 2021 5124 2699
rect 6900 2648 6920 5672
rect 6984 2648 7004 5672
rect 6900 2072 7004 2648
rect 3611 2020 6533 2021
rect 3611 -900 3612 2020
rect 6532 -900 6533 2020
rect 3611 -901 6533 -900
rect 2602 -1528 2706 -952
rect -687 -1580 2235 -1579
rect -687 -4500 -686 -1580
rect 2234 -4500 2235 -1580
rect -687 -4501 2235 -4500
rect -1696 -5128 -1592 -4552
rect -4985 -5180 -2063 -5179
rect -4985 -8100 -4984 -5180
rect -2064 -8100 -2063 -5180
rect -4985 -8101 -2063 -8100
rect -5994 -8300 -5890 -8152
rect -3576 -8300 -3472 -8101
rect -1696 -8152 -1676 -5128
rect -1612 -8152 -1592 -5128
rect 722 -5179 826 -4501
rect 2602 -4552 2622 -1528
rect 2686 -4552 2706 -1528
rect 5020 -1579 5124 -901
rect 6900 -952 6920 2072
rect 6984 -952 7004 2072
rect 6900 -1528 7004 -952
rect 3611 -1580 6533 -1579
rect 3611 -4500 3612 -1580
rect 6532 -4500 6533 -1580
rect 3611 -4501 6533 -4500
rect 2602 -5128 2706 -4552
rect -687 -5180 2235 -5179
rect -687 -8100 -686 -5180
rect 2234 -8100 2235 -5180
rect -687 -8101 2235 -8100
rect -1696 -8300 -1592 -8152
rect 722 -8300 826 -8101
rect 2602 -8152 2622 -5128
rect 2686 -8152 2706 -5128
rect 5020 -5179 5124 -4501
rect 6900 -4552 6920 -1528
rect 6984 -4552 7004 -1528
rect 6900 -5128 7004 -4552
rect 3611 -5180 6533 -5179
rect 3611 -8100 3612 -5180
rect 6532 -8100 6533 -5180
rect 3611 -8101 6533 -8100
rect 2602 -8300 2706 -8152
rect 5020 -8300 5124 -8101
rect 6900 -8152 6920 -5128
rect 6984 -8152 7004 -5128
rect 6900 -8300 7004 -8152
<< properties >>
string FIXED_BBOX 3732 5100 6812 8180
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 15.00 l 15.00 val 461.4 carea 2.00 cperi 0.19 nx 4 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
