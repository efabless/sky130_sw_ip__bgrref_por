magic
tech sky130A
timestamp 1717363523
<< pwell >>
rect -154 -1156 154 1156
<< mvnmos >>
rect -40 827 40 1027
rect -40 518 40 718
rect -40 209 40 409
rect -40 -100 40 100
rect -40 -409 40 -209
rect -40 -718 40 -518
rect -40 -1027 40 -827
<< mvndiff >>
rect -69 1021 -40 1027
rect -69 833 -63 1021
rect -46 833 -40 1021
rect -69 827 -40 833
rect 40 1021 69 1027
rect 40 833 46 1021
rect 63 833 69 1021
rect 40 827 69 833
rect -69 712 -40 718
rect -69 524 -63 712
rect -46 524 -40 712
rect -69 518 -40 524
rect 40 712 69 718
rect 40 524 46 712
rect 63 524 69 712
rect 40 518 69 524
rect -69 403 -40 409
rect -69 215 -63 403
rect -46 215 -40 403
rect -69 209 -40 215
rect 40 403 69 409
rect 40 215 46 403
rect 63 215 69 403
rect 40 209 69 215
rect -69 94 -40 100
rect -69 -94 -63 94
rect -46 -94 -40 94
rect -69 -100 -40 -94
rect 40 94 69 100
rect 40 -94 46 94
rect 63 -94 69 94
rect 40 -100 69 -94
rect -69 -215 -40 -209
rect -69 -403 -63 -215
rect -46 -403 -40 -215
rect -69 -409 -40 -403
rect 40 -215 69 -209
rect 40 -403 46 -215
rect 63 -403 69 -215
rect 40 -409 69 -403
rect -69 -524 -40 -518
rect -69 -712 -63 -524
rect -46 -712 -40 -524
rect -69 -718 -40 -712
rect 40 -524 69 -518
rect 40 -712 46 -524
rect 63 -712 69 -524
rect 40 -718 69 -712
rect -69 -833 -40 -827
rect -69 -1021 -63 -833
rect -46 -1021 -40 -833
rect -69 -1027 -40 -1021
rect 40 -833 69 -827
rect 40 -1021 46 -833
rect 63 -1021 69 -833
rect 40 -1027 69 -1021
<< mvndiffc >>
rect -63 833 -46 1021
rect 46 833 63 1021
rect -63 524 -46 712
rect 46 524 63 712
rect -63 215 -46 403
rect 46 215 63 403
rect -63 -94 -46 94
rect 46 -94 63 94
rect -63 -403 -46 -215
rect 46 -403 63 -215
rect -63 -712 -46 -524
rect 46 -712 63 -524
rect -63 -1021 -46 -833
rect 46 -1021 63 -833
<< mvpsubdiff >>
rect -136 1132 136 1138
rect -136 1115 -82 1132
rect 82 1115 136 1132
rect -136 1109 136 1115
rect -136 1084 -107 1109
rect -136 -1084 -130 1084
rect -113 -1084 -107 1084
rect 107 1084 136 1109
rect -136 -1109 -107 -1084
rect 107 -1084 113 1084
rect 130 -1084 136 1084
rect 107 -1109 136 -1084
rect -136 -1115 136 -1109
rect -136 -1132 -82 -1115
rect 82 -1132 136 -1115
rect -136 -1138 136 -1132
<< mvpsubdiffcont >>
rect -82 1115 82 1132
rect -130 -1084 -113 1084
rect 113 -1084 130 1084
rect -82 -1132 82 -1115
<< poly >>
rect -40 1063 40 1071
rect -40 1046 -32 1063
rect 32 1046 40 1063
rect -40 1027 40 1046
rect -40 808 40 827
rect -40 791 -32 808
rect 32 791 40 808
rect -40 783 40 791
rect -40 754 40 762
rect -40 737 -32 754
rect 32 737 40 754
rect -40 718 40 737
rect -40 499 40 518
rect -40 482 -32 499
rect 32 482 40 499
rect -40 474 40 482
rect -40 445 40 453
rect -40 428 -32 445
rect 32 428 40 445
rect -40 409 40 428
rect -40 190 40 209
rect -40 173 -32 190
rect 32 173 40 190
rect -40 165 40 173
rect -40 136 40 144
rect -40 119 -32 136
rect 32 119 40 136
rect -40 100 40 119
rect -40 -119 40 -100
rect -40 -136 -32 -119
rect 32 -136 40 -119
rect -40 -144 40 -136
rect -40 -173 40 -165
rect -40 -190 -32 -173
rect 32 -190 40 -173
rect -40 -209 40 -190
rect -40 -428 40 -409
rect -40 -445 -32 -428
rect 32 -445 40 -428
rect -40 -453 40 -445
rect -40 -482 40 -474
rect -40 -499 -32 -482
rect 32 -499 40 -482
rect -40 -518 40 -499
rect -40 -737 40 -718
rect -40 -754 -32 -737
rect 32 -754 40 -737
rect -40 -762 40 -754
rect -40 -791 40 -783
rect -40 -808 -32 -791
rect 32 -808 40 -791
rect -40 -827 40 -808
rect -40 -1046 40 -1027
rect -40 -1063 -32 -1046
rect 32 -1063 40 -1046
rect -40 -1071 40 -1063
<< polycont >>
rect -32 1046 32 1063
rect -32 791 32 808
rect -32 737 32 754
rect -32 482 32 499
rect -32 428 32 445
rect -32 173 32 190
rect -32 119 32 136
rect -32 -136 32 -119
rect -32 -190 32 -173
rect -32 -445 32 -428
rect -32 -499 32 -482
rect -32 -754 32 -737
rect -32 -808 32 -791
rect -32 -1063 32 -1046
<< locali >>
rect -130 1115 -82 1132
rect 82 1115 130 1132
rect -130 1084 -113 1115
rect 113 1084 130 1115
rect -40 1046 -32 1063
rect 32 1046 40 1063
rect -63 1021 -46 1029
rect -63 825 -46 833
rect 46 1021 63 1029
rect 46 825 63 833
rect -40 791 -32 808
rect 32 791 40 808
rect -40 737 -32 754
rect 32 737 40 754
rect -63 712 -46 720
rect -63 516 -46 524
rect 46 712 63 720
rect 46 516 63 524
rect -40 482 -32 499
rect 32 482 40 499
rect -40 428 -32 445
rect 32 428 40 445
rect -63 403 -46 411
rect -63 207 -46 215
rect 46 403 63 411
rect 46 207 63 215
rect -40 173 -32 190
rect 32 173 40 190
rect -40 119 -32 136
rect 32 119 40 136
rect -63 94 -46 102
rect -63 -102 -46 -94
rect 46 94 63 102
rect 46 -102 63 -94
rect -40 -136 -32 -119
rect 32 -136 40 -119
rect -40 -190 -32 -173
rect 32 -190 40 -173
rect -63 -215 -46 -207
rect -63 -411 -46 -403
rect 46 -215 63 -207
rect 46 -411 63 -403
rect -40 -445 -32 -428
rect 32 -445 40 -428
rect -40 -499 -32 -482
rect 32 -499 40 -482
rect -63 -524 -46 -516
rect -63 -720 -46 -712
rect 46 -524 63 -516
rect 46 -720 63 -712
rect -40 -754 -32 -737
rect 32 -754 40 -737
rect -40 -808 -32 -791
rect 32 -808 40 -791
rect -63 -833 -46 -825
rect -63 -1029 -46 -1021
rect 46 -833 63 -825
rect 46 -1029 63 -1021
rect -40 -1063 -32 -1046
rect 32 -1063 40 -1046
rect -130 -1115 -113 -1084
rect 113 -1115 130 -1084
rect -130 -1132 -82 -1115
rect 82 -1132 130 -1115
<< viali >>
rect -32 1046 32 1063
rect -63 833 -46 1021
rect 46 833 63 1021
rect -32 791 32 808
rect -32 737 32 754
rect -63 524 -46 712
rect 46 524 63 712
rect -32 482 32 499
rect -32 428 32 445
rect -63 215 -46 403
rect 46 215 63 403
rect -32 173 32 190
rect -32 119 32 136
rect -63 -94 -46 94
rect 46 -94 63 94
rect -32 -136 32 -119
rect -32 -190 32 -173
rect -63 -403 -46 -215
rect 46 -403 63 -215
rect -32 -445 32 -428
rect -32 -499 32 -482
rect -63 -712 -46 -524
rect 46 -712 63 -524
rect -32 -754 32 -737
rect -32 -808 32 -791
rect -63 -1021 -46 -833
rect 46 -1021 63 -833
rect -32 -1063 32 -1046
<< metal1 >>
rect -38 1063 38 1066
rect -38 1046 -32 1063
rect 32 1046 38 1063
rect -38 1043 38 1046
rect -66 1021 -43 1027
rect -66 833 -63 1021
rect -46 833 -43 1021
rect -66 827 -43 833
rect 43 1021 66 1027
rect 43 833 46 1021
rect 63 833 66 1021
rect 43 827 66 833
rect -38 808 38 811
rect -38 791 -32 808
rect 32 791 38 808
rect -38 788 38 791
rect -38 754 38 757
rect -38 737 -32 754
rect 32 737 38 754
rect -38 734 38 737
rect -66 712 -43 718
rect -66 524 -63 712
rect -46 524 -43 712
rect -66 518 -43 524
rect 43 712 66 718
rect 43 524 46 712
rect 63 524 66 712
rect 43 518 66 524
rect -38 499 38 502
rect -38 482 -32 499
rect 32 482 38 499
rect -38 479 38 482
rect -38 445 38 448
rect -38 428 -32 445
rect 32 428 38 445
rect -38 425 38 428
rect -66 403 -43 409
rect -66 215 -63 403
rect -46 215 -43 403
rect -66 209 -43 215
rect 43 403 66 409
rect 43 215 46 403
rect 63 215 66 403
rect 43 209 66 215
rect -38 190 38 193
rect -38 173 -32 190
rect 32 173 38 190
rect -38 170 38 173
rect -38 136 38 139
rect -38 119 -32 136
rect 32 119 38 136
rect -38 116 38 119
rect -66 94 -43 100
rect -66 -94 -63 94
rect -46 -94 -43 94
rect -66 -100 -43 -94
rect 43 94 66 100
rect 43 -94 46 94
rect 63 -94 66 94
rect 43 -100 66 -94
rect -38 -119 38 -116
rect -38 -136 -32 -119
rect 32 -136 38 -119
rect -38 -139 38 -136
rect -38 -173 38 -170
rect -38 -190 -32 -173
rect 32 -190 38 -173
rect -38 -193 38 -190
rect -66 -215 -43 -209
rect -66 -403 -63 -215
rect -46 -403 -43 -215
rect -66 -409 -43 -403
rect 43 -215 66 -209
rect 43 -403 46 -215
rect 63 -403 66 -215
rect 43 -409 66 -403
rect -38 -428 38 -425
rect -38 -445 -32 -428
rect 32 -445 38 -428
rect -38 -448 38 -445
rect -38 -482 38 -479
rect -38 -499 -32 -482
rect 32 -499 38 -482
rect -38 -502 38 -499
rect -66 -524 -43 -518
rect -66 -712 -63 -524
rect -46 -712 -43 -524
rect -66 -718 -43 -712
rect 43 -524 66 -518
rect 43 -712 46 -524
rect 63 -712 66 -524
rect 43 -718 66 -712
rect -38 -737 38 -734
rect -38 -754 -32 -737
rect 32 -754 38 -737
rect -38 -757 38 -754
rect -38 -791 38 -788
rect -38 -808 -32 -791
rect 32 -808 38 -791
rect -38 -811 38 -808
rect -66 -833 -43 -827
rect -66 -1021 -63 -833
rect -46 -1021 -43 -833
rect -66 -1027 -43 -1021
rect 43 -833 66 -827
rect 43 -1021 46 -833
rect 63 -1021 66 -833
rect 43 -1027 66 -1021
rect -38 -1046 38 -1043
rect -38 -1063 -32 -1046
rect 32 -1063 38 -1046
rect -38 -1066 38 -1063
<< properties >>
string FIXED_BBOX -121 -1123 121 1123
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2.0 l 0.8 m 7 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
