magic
tech sky130A
magscale 1 2
timestamp 1717613630
<< nwell >>
rect -672 -3780 -582 -2986
<< locali >>
rect 7082 -2491 10069 -2453
rect 10433 -2456 11133 -2453
rect 7082 -2551 7254 -2491
rect 10040 -2551 10069 -2491
rect 4856 -2620 4933 -2618
rect 4856 -2670 6961 -2620
rect 4856 -2726 4964 -2670
rect 6850 -2726 6961 -2670
rect -1971 -2769 -1764 -2766
rect -524 -2769 1782 -2768
rect -1971 -2863 1858 -2769
rect -1971 -3455 -1949 -2863
rect -1902 -2864 1858 -2863
rect -1902 -2934 -1812 -2864
rect 1696 -2934 1858 -2864
rect -1902 -3002 1858 -2934
rect -1902 -3084 -746 -3002
rect -1902 -3455 -1764 -3084
rect -1971 -3502 -1764 -3455
rect -1965 -4884 -1891 -3502
rect -783 -4884 -746 -3084
rect -1965 -4920 -746 -4884
rect -1965 -4974 -1854 -4920
rect -804 -4971 -746 -4920
rect -689 -3092 1858 -3002
rect -689 -3145 -362 -3092
rect -689 -3435 -466 -3145
rect -417 -3435 -362 -3145
rect -689 -3469 -362 -3435
rect 641 -3145 766 -3092
rect 641 -3435 662 -3145
rect 711 -3435 766 -3145
rect 641 -3465 766 -3435
rect -689 -3707 -471 -3469
rect 1762 -3707 1858 -3092
rect 1936 -2854 2998 -2835
rect 1936 -2903 2166 -2854
rect -689 -3710 -547 -3707
rect -689 -4971 -664 -3710
rect 1936 -4012 1971 -2903
rect 2026 -2926 2166 -2903
rect 2949 -2926 2998 -2854
rect 2026 -3046 2998 -2926
rect 2026 -4012 2079 -3046
rect 2860 -3137 2998 -3046
rect 2193 -3581 2435 -3145
rect 2525 -3581 2767 -3145
rect 1936 -4056 2079 -4012
rect -552 -4094 1344 -4056
rect -552 -4326 -528 -4094
rect -460 -4290 1344 -4094
rect -460 -4326 86 -4290
rect -552 -4380 86 -4326
rect -804 -4974 -664 -4971
rect -1965 -4994 -664 -4974
rect -1907 -5006 -664 -4994
rect -548 -5091 -436 -4380
rect -1984 -5134 -436 -5091
rect -1984 -5149 -592 -5134
rect -1984 -5500 -1922 -5149
rect -1983 -5522 -1922 -5500
rect -1866 -5507 -592 -5149
rect -536 -5334 -436 -5134
rect -536 -5472 -458 -5334
rect -186 -5472 62 -4380
rect 482 -4682 1344 -4290
rect 482 -5472 654 -4682
rect 1050 -4684 1344 -4682
rect 1050 -5404 1218 -4684
rect 1282 -5404 1344 -4684
rect 1050 -5472 1344 -5404
rect 1856 -4090 2079 -4056
rect 1856 -4114 2078 -4090
rect 1856 -5436 1898 -4114
rect 1960 -5436 2078 -4114
rect 2360 -5380 2602 -4944
rect 2860 -4946 2914 -3137
rect 2692 -5374 2914 -4946
rect 2970 -5374 2998 -3137
rect 4856 -2873 6961 -2726
rect 7082 -2759 10069 -2551
rect 7082 -2760 9091 -2759
rect 9222 -2760 10069 -2759
rect 10426 -2491 11133 -2456
rect 10426 -2551 10463 -2491
rect 11093 -2551 11133 -2491
rect 10426 -2760 11133 -2551
rect 4856 -4889 4933 -2873
rect 6881 -4138 6961 -2873
rect 7162 -3948 7251 -2760
rect 7538 -3729 7675 -2760
rect 7965 -3731 8102 -2760
rect 8391 -3332 8833 -2760
rect 9222 -3133 9481 -2760
rect 9819 -3133 10068 -2760
rect 8391 -3547 8698 -3332
rect 9222 -3449 9348 -3133
rect 9919 -3360 10068 -3133
rect 10426 -3136 10652 -2760
rect 10986 -3076 11132 -2760
rect 10985 -3129 11132 -3076
rect 10427 -3354 10527 -3136
rect 10985 -3345 11131 -3129
rect 9222 -3545 9408 -3449
rect 8391 -3725 8608 -3547
rect 8519 -3953 8608 -3725
rect 9669 -4119 9732 -4100
rect 6881 -4140 7353 -4138
rect 6881 -4192 7548 -4140
rect 5414 -4287 7548 -4192
rect 5424 -4889 5502 -4287
rect 6329 -4396 7548 -4287
rect 4856 -4973 5504 -4889
rect 4914 -4975 5504 -4973
rect 2692 -5382 2998 -5374
rect 1856 -5471 2078 -5436
rect 1734 -5472 2078 -5471
rect 2860 -5472 2998 -5382
rect -536 -5507 2998 -5472
rect -1866 -5522 2998 -5507
rect -1983 -5616 2998 -5522
rect -1983 -5682 -1931 -5616
rect 2904 -5682 2998 -5616
rect -1983 -5789 2998 -5682
rect -115 -5798 2998 -5789
rect 6329 -5537 6457 -4396
rect 7320 -5537 7548 -4396
rect 7940 -4198 8065 -4148
rect 7940 -5481 7999 -4198
rect 8037 -5481 8065 -4198
rect 7940 -5537 8065 -5481
rect 8468 -4198 8593 -4167
rect 8468 -5481 8526 -4198
rect 8564 -5481 8593 -4198
rect 8468 -5537 8593 -5481
rect 8600 -4374 8775 -4351
rect 8600 -5537 8911 -4374
rect 9205 -5537 9285 -4347
rect 9669 -4430 9679 -4119
rect 9722 -4239 9732 -4119
rect 9722 -4430 9838 -4239
rect 9669 -4446 9683 -4430
rect 9717 -4446 9732 -4430
rect 9383 -5537 9525 -4961
rect 9831 -5537 9973 -4958
rect 10296 -5537 10382 -4953
rect 6329 -5700 10382 -5537
rect 6329 -5748 6490 -5700
rect 10255 -5748 10382 -5700
rect -115 -5800 2890 -5798
rect 6329 -5799 10382 -5748
<< viali >>
rect 7254 -2551 10040 -2491
rect 4964 -2726 6850 -2670
rect -1949 -3455 -1902 -2863
rect -1812 -2934 1696 -2864
rect -1854 -4974 -804 -4920
rect -746 -4971 -689 -3002
rect -466 -3435 -417 -3145
rect 662 -3435 711 -3145
rect 1971 -4012 2026 -2903
rect 2166 -2926 2949 -2854
rect -528 -4326 -460 -4094
rect -1922 -5522 -1866 -5149
rect -592 -5507 -536 -5134
rect 1218 -5404 1282 -4684
rect 1898 -5436 1960 -4114
rect 2914 -5374 2970 -3137
rect 10463 -2551 11093 -2491
rect -1931 -5682 2904 -5616
rect 7999 -5481 8037 -4198
rect 8526 -5481 8564 -4198
rect 9679 -4430 9722 -4119
rect 6490 -5748 10255 -5700
<< metal1 >>
rect -1865 -2507 1863 -2466
rect -1865 -2710 -1803 -2507
rect 1801 -2533 1863 -2507
rect 1801 -2710 2029 -2533
rect 4114 -2641 4314 -2441
rect 4410 -2641 4610 -2441
rect 7082 -2491 10069 -2453
rect 10433 -2456 11133 -2453
rect 7082 -2511 7254 -2491
rect -1865 -2733 2029 -2710
rect -1865 -2766 1863 -2733
rect -1983 -2800 1863 -2766
rect -1983 -2863 1858 -2800
rect 4181 -2831 4250 -2641
rect 4481 -2835 4550 -2641
rect 4731 -2670 6895 -2620
rect 4731 -2726 4964 -2670
rect 6850 -2726 6895 -2670
rect -1983 -3455 -1949 -2863
rect -1902 -2864 1858 -2863
rect -1902 -2934 -1812 -2864
rect 1696 -2934 1858 -2864
rect -1902 -3002 1858 -2934
rect -1902 -3084 -746 -3002
rect -1902 -3455 -1764 -3084
rect -1983 -3502 -1764 -3455
rect -1983 -4886 -1906 -3502
rect -1398 -3521 -1303 -3218
rect -904 -3521 -836 -3286
rect -1718 -3574 -836 -3521
rect -1844 -4126 -1776 -3890
rect -1398 -4126 -1303 -3815
rect -904 -4079 -836 -3574
rect -1844 -4179 -942 -4126
rect -1844 -4683 -1776 -4179
rect -1393 -4735 -1298 -4419
rect -936 -4735 -855 -4731
rect -1723 -4788 -855 -4735
rect -936 -4789 -855 -4788
rect -773 -4886 -746 -3084
rect -1983 -4920 -746 -4886
rect -1983 -4974 -1854 -4920
rect -804 -4971 -746 -4920
rect -689 -3092 1858 -3002
rect -689 -3145 -362 -3092
rect -689 -3435 -466 -3145
rect -417 -3435 -362 -3145
rect 641 -3145 766 -3092
rect -689 -3469 -362 -3435
rect -689 -3707 -471 -3469
rect -689 -3710 -547 -3707
rect -689 -4971 -662 -3710
rect 30 -3832 136 -3208
rect 516 -3660 588 -3282
rect 641 -3435 662 -3145
rect 711 -3435 766 -3145
rect 641 -3465 766 -3435
rect 516 -3732 788 -3660
rect 27 -3928 431 -3832
rect -420 -4006 298 -3968
rect -804 -4974 -662 -4971
rect -1983 -5004 -662 -4974
rect -1915 -5005 -662 -5004
rect -773 -5008 -662 -5005
rect -548 -4094 -436 -4056
rect -548 -4326 -528 -4094
rect -460 -4326 -436 -4094
rect -548 -5091 -436 -4326
rect -376 -4449 -200 -4448
rect -376 -4490 -191 -4449
rect -1984 -5134 -436 -5091
rect -1984 -5149 -592 -5134
rect -1984 -5500 -1922 -5149
rect -1983 -5522 -1922 -5500
rect -1866 -5507 -592 -5149
rect -536 -5330 -436 -5134
rect -536 -5472 -458 -5330
rect -233 -5368 -191 -4490
rect -394 -5410 -186 -5368
rect 126 -5393 198 -4482
rect 260 -5348 298 -4006
rect 358 -5278 430 -3928
rect 716 -5395 788 -3732
rect 1146 -3832 1252 -3214
rect 1634 -3658 1702 -3292
rect 1398 -3726 1702 -3658
rect 1762 -3707 1858 -3092
rect 1936 -2854 2998 -2835
rect 1936 -2903 2166 -2854
rect 1398 -3832 1466 -3726
rect 1146 -3918 1467 -3832
rect 1146 -3920 1252 -3918
rect 1050 -4684 1300 -4628
rect 890 -5331 932 -4841
rect 1050 -5404 1218 -4684
rect 1282 -5404 1300 -4684
rect 1398 -5278 1466 -3918
rect 1936 -4012 1971 -2903
rect 2026 -2926 2166 -2903
rect 2949 -2926 2998 -2854
rect 2026 -2928 2998 -2926
rect 4731 -2873 6895 -2726
rect 7082 -2697 7151 -2511
rect 10040 -2551 10069 -2491
rect 9985 -2697 10069 -2551
rect 7082 -2759 10069 -2697
rect 7082 -2760 9091 -2759
rect 9339 -2760 10069 -2759
rect 10426 -2491 11133 -2456
rect 10426 -2551 10463 -2491
rect 11093 -2551 11133 -2491
rect 10426 -2760 11133 -2551
rect 4731 -2928 4940 -2873
rect 2026 -3046 4940 -2928
rect 2026 -4012 2079 -3046
rect 2860 -3137 4940 -3046
rect 2193 -3581 2435 -3145
rect 2525 -3581 2767 -3145
rect 1936 -4057 2079 -4012
rect 1932 -4058 2079 -4057
rect 1856 -4090 2079 -4058
rect 1856 -4114 2075 -4090
rect 1580 -5331 1618 -4202
rect 1726 -5280 1783 -4262
rect 1050 -5472 1300 -5404
rect 1856 -5436 1898 -4114
rect 1960 -5436 2075 -4114
rect 2360 -5380 2602 -4944
rect 2860 -4946 2914 -3137
rect 2692 -5374 2914 -4946
rect 2970 -5374 3113 -3137
rect 5147 -4085 5190 -2943
rect 5358 -3060 5468 -3044
rect 5358 -3666 5468 -3199
rect 5147 -4099 5195 -4085
rect 4858 -4370 4967 -4355
rect 4628 -4853 4814 -4818
rect 4779 -5328 4814 -4853
rect 4858 -5154 4967 -4508
rect 5151 -4805 5195 -4099
rect 5358 -4578 5468 -3805
rect 5639 -4101 5682 -2945
rect 5853 -3259 5960 -3241
rect 5853 -3887 5960 -3398
rect 5358 -4724 5468 -4717
rect 5853 -4974 5960 -4026
rect 6126 -4106 6169 -2950
rect 6330 -3060 6440 -3044
rect 6330 -3666 6440 -3199
rect 6330 -4578 6440 -3805
rect 6608 -4106 6651 -2950
rect 7082 -3877 7129 -2760
rect 7322 -3964 7371 -2937
rect 7440 -3791 7469 -2863
rect 7538 -3729 7675 -2760
rect 7747 -3710 7796 -2932
rect 7747 -3791 7803 -3710
rect 7866 -3791 7895 -2863
rect 7965 -3731 8102 -2760
rect 7411 -3834 7931 -3791
rect 7083 -4013 7371 -3964
rect 7083 -4272 7129 -4013
rect 7751 -4063 7802 -3834
rect 8163 -3980 8228 -2930
rect 8288 -3798 8319 -2857
rect 8391 -3725 8528 -2760
rect 8658 -3332 8833 -2760
rect 8950 -3371 9001 -2863
rect 9114 -3371 9158 -2939
rect 9339 -3133 9481 -2760
rect 9551 -3197 9585 -2875
rect 9710 -3197 9744 -2878
rect 9819 -3133 10068 -2760
rect 10426 -3136 10652 -2760
rect 10724 -3189 10758 -2877
rect 10889 -3183 10923 -2878
rect 10986 -3129 11132 -2760
rect 10769 -3189 10923 -3183
rect 10185 -3193 10923 -3189
rect 8879 -3418 9158 -3371
rect 8879 -3420 8886 -3418
rect 9030 -3420 9158 -3418
rect 9114 -3683 9158 -3420
rect 9537 -3230 9757 -3197
rect 10185 -3222 10928 -3193
rect 9537 -3598 9570 -3230
rect 10185 -3492 10218 -3222
rect 10724 -3225 10928 -3222
rect 10769 -3226 10928 -3225
rect 10769 -3228 10918 -3226
rect 9626 -3540 10218 -3492
rect 9537 -3631 10073 -3598
rect 9114 -3729 9821 -3683
rect 6755 -4318 7129 -4272
rect 7183 -4114 7802 -4063
rect 8145 -3997 8228 -3980
rect 8145 -4058 9015 -3997
rect 6330 -4724 6440 -4717
rect 5853 -5137 5960 -5120
rect 4858 -5283 4967 -5266
rect 5211 -5328 5246 -5246
rect 4779 -5363 5246 -5328
rect 2692 -5382 3113 -5374
rect 1856 -5471 2075 -5436
rect 1734 -5472 2075 -5471
rect 2860 -5472 3113 -5382
rect 6656 -5409 6685 -4501
rect 6755 -5362 6801 -4318
rect 7082 -5409 7111 -4506
rect 7183 -5366 7234 -4114
rect 7401 -5409 7443 -4145
rect 7940 -4198 8065 -4148
rect 7614 -5355 7668 -4359
rect 6656 -5445 7443 -5409
rect 7782 -5429 7824 -4283
rect 6658 -5451 7443 -5445
rect -536 -5507 3113 -5472
rect -1866 -5522 3113 -5507
rect -1983 -5530 3113 -5522
rect 7940 -5481 7999 -4198
rect 8037 -5481 8065 -4198
rect 8145 -5357 8199 -4058
rect 8468 -4198 8593 -4167
rect 8305 -5427 8347 -4281
rect -1983 -5537 6597 -5530
rect 7940 -5537 8065 -5481
rect 8468 -5481 8526 -4198
rect 8564 -5481 8593 -4198
rect 8468 -5537 8593 -5481
rect 8769 -5537 8911 -4374
rect 8978 -4488 9015 -4058
rect 9669 -4119 9732 -4100
rect 9669 -4430 9679 -4119
rect 9722 -4239 9732 -4119
rect 9775 -4239 9821 -3729
rect 9722 -4430 9838 -4239
rect 9669 -4446 9732 -4430
rect 9893 -4488 9930 -4157
rect 10040 -4238 10073 -3631
rect 8978 -4524 9953 -4488
rect 8978 -5425 9015 -4524
rect 9992 -4627 10073 -4238
rect 9072 -4722 10073 -4627
rect 9072 -5366 9137 -4722
rect 10040 -4765 10073 -4722
rect 9601 -4798 10073 -4765
rect 9383 -5537 9525 -4961
rect 9601 -5430 9634 -4798
rect 10144 -4840 10218 -3540
rect 9711 -4888 10218 -4840
rect 9711 -5360 9759 -4888
rect 10185 -4947 10218 -4888
rect 9831 -5537 9973 -4958
rect 10051 -4980 10218 -4947
rect 10300 -3939 10348 -3558
rect 10555 -3939 10755 -3885
rect 10300 -4048 10755 -3939
rect 10051 -5432 10084 -4980
rect 10300 -5018 10348 -4048
rect 10555 -4085 10755 -4048
rect 10144 -5066 10348 -5018
rect 10144 -5365 10192 -5066
rect -1983 -5616 10309 -5537
rect -1983 -5682 -1931 -5616
rect 2904 -5682 10309 -5616
rect -1983 -5700 10309 -5682
rect -1983 -5748 6490 -5700
rect 10255 -5748 10309 -5700
rect -1983 -5772 10309 -5748
rect -116 -5789 10309 -5772
rect -115 -5799 10309 -5789
rect -115 -5800 6597 -5799
rect 2823 -5804 6597 -5800
<< via1 >>
rect -1803 -2710 1801 -2507
rect 7151 -2551 7254 -2511
rect 7254 -2551 9985 -2511
rect 7151 -2697 9985 -2551
rect 3307 -3890 4604 -3762
rect 5358 -3199 5468 -3060
rect 5358 -3805 5468 -3666
rect 4858 -4508 4967 -4370
rect 5853 -3398 5960 -3259
rect 5853 -4026 5960 -3887
rect 5358 -4717 5468 -4578
rect 6330 -3199 6440 -3060
rect 6330 -3805 6440 -3666
rect 6330 -4717 6440 -4578
rect 5853 -5120 5960 -4974
rect 4858 -5266 4967 -5154
<< metal2 >>
rect -1879 -2507 10067 -2441
rect -1879 -2710 -1803 -2507
rect 1801 -2511 10067 -2507
rect 1801 -2697 7151 -2511
rect 9985 -2697 10067 -2511
rect 1801 -2710 10067 -2697
rect -1879 -2751 10067 -2710
rect 3562 -3709 3937 -2751
rect 4187 -3537 4245 -2838
rect 4492 -3438 4536 -2833
rect 4980 -3199 5358 -3060
rect 5468 -3199 6330 -3060
rect 6440 -3199 6448 -3060
rect 6522 -3199 7010 -3060
rect 4980 -3398 5853 -3259
rect 5960 -3398 6808 -3259
rect 4492 -3482 6420 -3438
rect 4187 -3595 6270 -3537
rect 6376 -3540 6420 -3482
rect 6376 -3584 6595 -3540
rect 6870 -3666 7009 -3199
rect 9611 -3541 9675 -2981
rect 10779 -3470 10843 -2974
rect 10300 -3534 10843 -3470
rect 3225 -3762 4690 -3709
rect 26 -3922 1469 -3833
rect 3225 -3890 3307 -3762
rect 4604 -3890 4690 -3762
rect 4982 -3805 5358 -3666
rect 5468 -3805 6330 -3666
rect 6440 -3805 6450 -3666
rect 6521 -3805 7009 -3666
rect -328 -3923 -258 -3922
rect -441 -4019 -118 -3923
rect 3225 -3981 4690 -3890
rect -328 -4567 -258 -4019
rect 4986 -4026 5853 -3887
rect 5960 -4026 6814 -3887
rect 4628 -4228 5694 -4137
rect 4546 -4274 5694 -4228
rect 4546 -4365 4765 -4274
rect -888 -4722 -255 -4567
rect 4557 -4580 4751 -4464
rect 4842 -4508 4858 -4370
rect 4967 -4508 5393 -4370
rect 5557 -4578 5694 -4274
rect 6456 -4578 6595 -4577
rect -330 -4864 -255 -4722
rect 1724 -5235 2256 -4962
rect 3146 -5154 3258 -4788
rect 4635 -4974 4751 -4580
rect 5005 -4717 5358 -4578
rect 5468 -4717 6330 -4578
rect 6440 -4717 6596 -4578
rect 6456 -4860 6595 -4717
rect 6870 -4859 7009 -3805
rect 7070 -3999 7142 -3746
rect 7290 -3849 8414 -3782
rect 7070 -4071 7453 -3999
rect 7381 -4277 7453 -4071
rect 8138 -4511 8489 -4365
rect 4635 -5106 5853 -4974
rect 4638 -5120 5853 -5106
rect 5960 -5120 7980 -4974
rect 3146 -5266 4858 -5154
rect 4967 -5266 4980 -5154
rect 5296 -5226 9114 -5221
rect 5326 -5276 9114 -5226
rect -230 -5321 3139 -5315
rect -230 -5382 4749 -5321
rect -230 -5393 3139 -5382
rect 4688 -5397 4749 -5382
rect 4688 -5458 8422 -5397
use por_via_2cut  por_via_2cut_0
timestamp 1717613630
transform 0 1 12943 -1 0 12197
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_1
timestamp 1717613630
transform 0 1 14397 -1 0 12197
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_2
timestamp 1717613630
transform -1 0 20668 0 -1 -10745
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_3
timestamp 1717613630
transform 0 1 13917 -1 0 12200
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_4
timestamp 1717613630
transform 0 1 13204 -1 0 12420
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_5
timestamp 1717613630
transform 0 1 14659 -1 0 12416
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_6
timestamp 1717613630
transform 0 1 14171 -1 0 12418
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_7
timestamp 1717613630
transform 0 1 13686 -1 0 12413
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_8
timestamp 1717613630
transform 0 1 13197 -1 0 13028
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_9
timestamp 1717613630
transform 0 1 12941 -1 0 12829
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_10
timestamp 1717613630
transform 0 1 13686 -1 0 13026
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_11
timestamp 1717613630
transform 0 1 13426 -1 0 12825
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_12
timestamp 1717613630
transform 0 1 14402 -1 0 12824
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_13
timestamp 1717613630
transform 0 1 13915 -1 0 12823
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_14
timestamp 1717613630
transform 0 1 14175 -1 0 13020
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_15
timestamp 1717613630
transform 0 1 13195 -1 0 11717
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_16
timestamp 1717613630
transform 0 1 14659 -1 0 13024
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_17
timestamp 1717613630
transform 0 1 12943 -1 0 11505
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_18
timestamp 1717613630
transform 0 1 15320 -1 0 11946
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_19
timestamp 1717613630
transform 0 1 15210 -1 0 12354
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_20
timestamp 1717613630
transform 0 1 15006 -1 0 12338
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_21
timestamp 1717613630
transform -1 0 21420 0 -1 -13152
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_22
timestamp 1717613630
transform 0 1 17543 -1 0 12681
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_23
timestamp 1717613630
transform 0 1 17545 -1 0 13110
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_24
timestamp 1717613630
transform 0 1 18723 -1 0 13103
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_25
timestamp 1717613630
transform 0 1 18230 -1 0 12648
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_26
timestamp 1717613630
transform -1 0 24499 0 -1 -11716
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_27
timestamp 1717613630
transform 0 1 13429 -1 0 12199
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_28
timestamp 1717613630
transform -1 0 20373 0 -1 -10747
box 16088 -7932 16222 -7868
use por_via_4cut  por_via_4cut_0
timestamp 1717613630
transform 0 1 8061 -1 0 10839
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_1
timestamp 1717613630
transform 0 1 7019 -1 0 11490
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_2
timestamp 1717613630
transform -1 0 15801 0 -1 -11868
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_3
timestamp 1717613630
transform -1 0 16958 0 -1 -13253
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_4
timestamp 1717613630
transform 0 -1 -5679 1 0 -21185
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_5
timestamp 1717613630
transform -1 0 16264 0 -1 -11776
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_6
timestamp 1717613630
transform -1 0 17631 0 -1 -13253
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_7
timestamp 1717613630
transform 0 -1 -6136 1 0 -21185
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_8
timestamp 1717613630
transform -1 0 21256 0 -1 -11471
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_9
timestamp 1717613630
transform -1 0 22713 0 -1 -11465
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_10
timestamp 1717613630
transform -1 0 21753 0 -1 -11467
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_11
timestamp 1717613630
transform -1 0 22223 0 -1 -11469
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_12
timestamp 1717613630
transform 0 -1 -1337 1 0 -20823
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_13
timestamp 1717613630
transform 0 -1 -260 1 0 -21067
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_14
timestamp 1717613630
transform 0 -1 1202 1 0 -21226
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_15
timestamp 1717613630
transform 0 -1 -903 1 0 -20819
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_16
timestamp 1717613630
transform 0 1 7702 -1 0 10833
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_17
timestamp 1717613630
transform -1 0 17397 0 -1 -11776
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_18
timestamp 1717613630
transform -1 0 23858 0 -1 -13324
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_19
timestamp 1717613630
transform -1 0 24358 0 -1 -13328
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_20
timestamp 1717613630
transform 0 -1 269 1 0 -20579
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_21
timestamp 1717613630
transform 0 1 7608 -1 0 11375
box 15948 -7932 16222 -7868
use sky130_fd_pr__nfet_01v8_B8TQK3  sky130_fd_pr__nfet_01v8_B8TQK3_0 paramcells
timestamp 1717527227
transform -1 0 5176 0 1 -3526
box -296 -719 296 719
use sky130_fd_pr__nfet_01v8_B8TQK3  sky130_fd_pr__nfet_01v8_B8TQK3_1
timestamp 1717527227
transform -1 0 6148 0 1 -3526
box -296 -719 296 719
use sky130_fd_pr__nfet_01v8_B8TQK3  sky130_fd_pr__nfet_01v8_B8TQK3_2
timestamp 1717527227
transform -1 0 5662 0 1 -3526
box -296 -719 296 719
use mux2to1  x1
timestamp 1717613630
transform -1 0 5102 0 1 -4041
box 404 -1761 1956 334
use sky130_fd_pr__nfet_g5v0d10v5_T4TNG7  XM1 paramcells
timestamp 1717613630
transform -1 0 7798 0 1 -4856
box -333 -767 338 767
use sky130_fd_pr__pfet_g5v0d10v5_KL3SY6  XM2 paramcells
timestamp 1717527227
transform -1 0 7454 0 1 -3328
box -308 -697 308 697
use sky130_fd_pr__pfet_g5v0d10v5_KL3SY6  XM3
timestamp 1717527227
transform -1 0 7880 0 1 -3328
box -308 -697 308 697
use sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3  XM4 paramcells
timestamp 1717613630
transform 1 0 7103 0 1 -4978
box -283 -658 283 658
use sky130_fd_pr__pfet_g5v0d10v5_VHBZVD  XM5 paramcells
timestamp 1717613630
transform 1 0 -1330 0 1 -3383
box -658 -397 658 397
use sky130_fd_pr__nfet_g5v0d10v5_T4TNG7  XM6
timestamp 1717613630
transform 1 0 8334 0 1 -4856
box -333 -767 338 767
use sky130_fd_pr__pfet_g5v0d10v5_KL3SY6  XM7
timestamp 1717527227
transform 1 0 8306 0 1 -3328
box -308 -697 308 697
use sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3  XM8
timestamp 1717613630
transform 1 0 6667 0 1 -4978
box -283 -658 283 658
use sky130_fd_pr__nfet_01v8_QGMAL3  XM9 paramcells
timestamp 1717527227
transform 1 0 5176 0 1 -4549
box -296 -410 296 410
use sky130_fd_pr__nfet_01v8_B8TQK3  XM10
timestamp 1717527227
transform 1 0 6634 0 1 -3526
box -296 -719 296 719
use sky130_fd_pr__pfet_g5v0d10v5_VHBZVD  XM11
timestamp 1717613630
transform 1 0 -1330 0 1 -3987
box -658 -397 658 397
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM12 paramcells
timestamp 1717613630
transform 1 0 9619 0 1 -5270
box -288 -358 288 358
use sky130_fd_pr__pfet_g5v0d10v5_KLNSY6  XM13 paramcells
timestamp 1717527227
transform 1 0 9647 0 1 -3042
box -387 -397 387 397
use sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3  XM14
timestamp 1717613630
transform 1 0 8998 0 1 -4967
box -283 -658 283 658
use sky130_fd_pr__pfet_g5v0d10v5_KLAZY6  XM15 paramcells
timestamp 1717527227
transform 1 0 9913 0 1 -4338
box -308 -397 308 397
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM16
timestamp 1717613630
transform 1 0 10065 0 1 -5270
box -288 -358 288 358
use sky130_fd_pr__pfet_g5v0d10v5_KLNSY6  XM17
timestamp 1717527227
transform 1 0 10821 0 1 -3042
box -387 -397 387 397
use sky130_fd_pr__pfet_g5v0d10v5_FGK6VM  XM19 paramcells
timestamp 1717527227
transform 1 0 8971 0 1 -3136
box -358 -497 358 497
use sky130_fd_pr__pfet_g5v0d10v5_VHBZVD  XM20
timestamp 1717613630
transform 1 0 -1330 0 1 -4591
box -658 -397 658 397
use sky130_fd_pr__pfet_g5v0d10v5_VHBZVD  XM23
timestamp 1717613630
transform 1 0 1202 0 1 -3383
box -658 -397 658 397
use sky130_fd_pr__pfet_g5v0d10v5_VHBZVD  XM24
timestamp 1717613630
transform 1 0 76 0 1 -3383
box -658 -397 658 397
use sky130_fd_pr__nfet_g5v0d10v5_YYAQG7  XM25 paramcells
timestamp 1717613630
transform 1 0 914 0 1 -5082
box -328 -458 328 458
use sky130_fd_pr__nfet_g5v0d10v5_T4TNG7  XM26
timestamp 1717613630
transform 1 0 1600 0 1 -4773
box -333 -767 338 767
use sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3  XM27
timestamp 1717613630
transform 1 0 280 0 1 -4884
box -283 -658 283 658
use sky130_fd_pr__nfet_01v8_SALWK2  XM28 paramcells
timestamp 1717613630
transform 1 0 -364 0 1 -4930
box -226 -610 226 610
use sky130_fd_pr__res_xhigh_po_0p35_FVGVKR  XR12 paramcells
timestamp 1717613630
transform 1 0 2478 0 1 -4264
box -450 -1282 450 1282
<< labels >>
flabel metal2 4836 -3570 4836 -3570 0 FreeSans 400 0 0 0 Vinn
flabel metal2 4833 -3461 4833 -3461 0 FreeSans 400 0 0 0 Vinp
flabel via1 4863 -4442 4863 -4442 0 FreeSans 400 0 0 0 VY
flabel metal2 5605 -4649 5605 -4649 0 FreeSans 400 0 0 0 VD
flabel metal2 5880 -5436 5880 -5436 0 FreeSans 400 0 0 0 vbn
flabel metal1 8630 -4027 8630 -4027 0 FreeSans 400 0 0 0 vo
flabel metal2 6195 -5048 6195 -5048 0 FreeSans 400 0 0 0 VS
flabel metal2 8000 -3820 8000 -3820 0 FreeSans 400 0 0 0 vt
flabel via1 8651 -2599 8651 -2599 0 FreeSans 400 0 0 0 AVDD
flabel metal1 614 -2821 614 -2821 0 FreeSans 400 0 0 0 AVDD
flabel metal1 941 -5695 941 -5695 0 FreeSans 400 0 0 0 VSS
flabel metal2 3096 -5356 3096 -5356 0 FreeSans 400 0 0 0 vbn
flabel metal1 1829 -2733 2029 -2533 0 FreeSans 256 0 0 0 AVDD
port 4 nsew
flabel metal1 4821 -5777 5021 -5577 0 FreeSans 256 0 0 0 VSS
port 3 nsew
flabel metal1 10555 -4085 10755 -3885 0 FreeSans 256 0 0 0 RST
port 2 nsew
flabel metal1 4114 -2641 4314 -2441 0 FreeSans 256 0 0 0 Vinn
port 0 nsew
flabel metal1 4410 -2641 4610 -2441 0 FreeSans 256 0 0 0 Vinp
port 1 nsew
flabel metal1 8345 -5667 8345 -5667 0 FreeSans 400 0 0 0 VSS
flabel metal1 5623 -2770 5623 -2770 0 FreeSans 400 0 0 0 VSS
flabel metal1 10494 -3992 10494 -3992 0 FreeSans 400 0 0 0 RST
flabel metal1 9420 -4671 9420 -4671 0 FreeSans 400 0 0 0 vo1
flabel metal1 10893 -2737 11093 -2537 0 FreeSans 256 0 0 0 DVDD
port 5 nsew
flabel metal1 10776 -2599 10776 -2599 0 FreeSans 400 0 0 0 DVDD
<< end >>
