magic
tech sky130A
magscale 1 2
timestamp 1717443058
<< error_p >>
rect -2477 151 -2419 157
rect -2285 151 -2227 157
rect -2093 151 -2035 157
rect -1901 151 -1843 157
rect -1709 151 -1651 157
rect -1517 151 -1459 157
rect -1325 151 -1267 157
rect -1133 151 -1075 157
rect -941 151 -883 157
rect -749 151 -691 157
rect -557 151 -499 157
rect -365 151 -307 157
rect -173 151 -115 157
rect 19 151 77 157
rect 211 151 269 157
rect 403 151 461 157
rect 595 151 653 157
rect 787 151 845 157
rect 979 151 1037 157
rect 1171 151 1229 157
rect 1363 151 1421 157
rect 1555 151 1613 157
rect 1747 151 1805 157
rect 1939 151 1997 157
rect 2131 151 2189 157
rect 2323 151 2381 157
rect 2515 151 2573 157
rect -2477 117 -2465 151
rect -2285 117 -2273 151
rect -2093 117 -2081 151
rect -1901 117 -1889 151
rect -1709 117 -1697 151
rect -1517 117 -1505 151
rect -1325 117 -1313 151
rect -1133 117 -1121 151
rect -941 117 -929 151
rect -749 117 -737 151
rect -557 117 -545 151
rect -365 117 -353 151
rect -173 117 -161 151
rect 19 117 31 151
rect 211 117 223 151
rect 403 117 415 151
rect 595 117 607 151
rect 787 117 799 151
rect 979 117 991 151
rect 1171 117 1183 151
rect 1363 117 1375 151
rect 1555 117 1567 151
rect 1747 117 1759 151
rect 1939 117 1951 151
rect 2131 117 2143 151
rect 2323 117 2335 151
rect 2515 117 2527 151
rect -2477 111 -2419 117
rect -2285 111 -2227 117
rect -2093 111 -2035 117
rect -1901 111 -1843 117
rect -1709 111 -1651 117
rect -1517 111 -1459 117
rect -1325 111 -1267 117
rect -1133 111 -1075 117
rect -941 111 -883 117
rect -749 111 -691 117
rect -557 111 -499 117
rect -365 111 -307 117
rect -173 111 -115 117
rect 19 111 77 117
rect 211 111 269 117
rect 403 111 461 117
rect 595 111 653 117
rect 787 111 845 117
rect 979 111 1037 117
rect 1171 111 1229 117
rect 1363 111 1421 117
rect 1555 111 1613 117
rect 1747 111 1805 117
rect 1939 111 1997 117
rect 2131 111 2189 117
rect 2323 111 2381 117
rect 2515 111 2573 117
rect -2573 -117 -2515 -111
rect -2381 -117 -2323 -111
rect -2189 -117 -2131 -111
rect -1997 -117 -1939 -111
rect -1805 -117 -1747 -111
rect -1613 -117 -1555 -111
rect -1421 -117 -1363 -111
rect -1229 -117 -1171 -111
rect -1037 -117 -979 -111
rect -845 -117 -787 -111
rect -653 -117 -595 -111
rect -461 -117 -403 -111
rect -269 -117 -211 -111
rect -77 -117 -19 -111
rect 115 -117 173 -111
rect 307 -117 365 -111
rect 499 -117 557 -111
rect 691 -117 749 -111
rect 883 -117 941 -111
rect 1075 -117 1133 -111
rect 1267 -117 1325 -111
rect 1459 -117 1517 -111
rect 1651 -117 1709 -111
rect 1843 -117 1901 -111
rect 2035 -117 2093 -111
rect 2227 -117 2285 -111
rect 2419 -117 2477 -111
rect -2573 -151 -2561 -117
rect -2381 -151 -2369 -117
rect -2189 -151 -2177 -117
rect -1997 -151 -1985 -117
rect -1805 -151 -1793 -117
rect -1613 -151 -1601 -117
rect -1421 -151 -1409 -117
rect -1229 -151 -1217 -117
rect -1037 -151 -1025 -117
rect -845 -151 -833 -117
rect -653 -151 -641 -117
rect -461 -151 -449 -117
rect -269 -151 -257 -117
rect -77 -151 -65 -117
rect 115 -151 127 -117
rect 307 -151 319 -117
rect 499 -151 511 -117
rect 691 -151 703 -117
rect 883 -151 895 -117
rect 1075 -151 1087 -117
rect 1267 -151 1279 -117
rect 1459 -151 1471 -117
rect 1651 -151 1663 -117
rect 1843 -151 1855 -117
rect 2035 -151 2047 -117
rect 2227 -151 2239 -117
rect 2419 -151 2431 -117
rect -2573 -157 -2515 -151
rect -2381 -157 -2323 -151
rect -2189 -157 -2131 -151
rect -1997 -157 -1939 -151
rect -1805 -157 -1747 -151
rect -1613 -157 -1555 -151
rect -1421 -157 -1363 -151
rect -1229 -157 -1171 -151
rect -1037 -157 -979 -151
rect -845 -157 -787 -151
rect -653 -157 -595 -151
rect -461 -157 -403 -151
rect -269 -157 -211 -151
rect -77 -157 -19 -151
rect 115 -157 173 -151
rect 307 -157 365 -151
rect 499 -157 557 -151
rect 691 -157 749 -151
rect 883 -157 941 -151
rect 1075 -157 1133 -151
rect 1267 -157 1325 -151
rect 1459 -157 1517 -151
rect 1651 -157 1709 -151
rect 1843 -157 1901 -151
rect 2035 -157 2093 -151
rect 2227 -157 2285 -151
rect 2419 -157 2477 -151
<< nwell >>
rect -2759 -289 2759 289
<< pmos >>
rect -2559 -70 -2529 70
rect -2463 -70 -2433 70
rect -2367 -70 -2337 70
rect -2271 -70 -2241 70
rect -2175 -70 -2145 70
rect -2079 -70 -2049 70
rect -1983 -70 -1953 70
rect -1887 -70 -1857 70
rect -1791 -70 -1761 70
rect -1695 -70 -1665 70
rect -1599 -70 -1569 70
rect -1503 -70 -1473 70
rect -1407 -70 -1377 70
rect -1311 -70 -1281 70
rect -1215 -70 -1185 70
rect -1119 -70 -1089 70
rect -1023 -70 -993 70
rect -927 -70 -897 70
rect -831 -70 -801 70
rect -735 -70 -705 70
rect -639 -70 -609 70
rect -543 -70 -513 70
rect -447 -70 -417 70
rect -351 -70 -321 70
rect -255 -70 -225 70
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
rect 225 -70 255 70
rect 321 -70 351 70
rect 417 -70 447 70
rect 513 -70 543 70
rect 609 -70 639 70
rect 705 -70 735 70
rect 801 -70 831 70
rect 897 -70 927 70
rect 993 -70 1023 70
rect 1089 -70 1119 70
rect 1185 -70 1215 70
rect 1281 -70 1311 70
rect 1377 -70 1407 70
rect 1473 -70 1503 70
rect 1569 -70 1599 70
rect 1665 -70 1695 70
rect 1761 -70 1791 70
rect 1857 -70 1887 70
rect 1953 -70 1983 70
rect 2049 -70 2079 70
rect 2145 -70 2175 70
rect 2241 -70 2271 70
rect 2337 -70 2367 70
rect 2433 -70 2463 70
rect 2529 -70 2559 70
<< pdiff >>
rect -2621 58 -2559 70
rect -2621 -58 -2609 58
rect -2575 -58 -2559 58
rect -2621 -70 -2559 -58
rect -2529 58 -2463 70
rect -2529 -58 -2513 58
rect -2479 -58 -2463 58
rect -2529 -70 -2463 -58
rect -2433 58 -2367 70
rect -2433 -58 -2417 58
rect -2383 -58 -2367 58
rect -2433 -70 -2367 -58
rect -2337 58 -2271 70
rect -2337 -58 -2321 58
rect -2287 -58 -2271 58
rect -2337 -70 -2271 -58
rect -2241 58 -2175 70
rect -2241 -58 -2225 58
rect -2191 -58 -2175 58
rect -2241 -70 -2175 -58
rect -2145 58 -2079 70
rect -2145 -58 -2129 58
rect -2095 -58 -2079 58
rect -2145 -70 -2079 -58
rect -2049 58 -1983 70
rect -2049 -58 -2033 58
rect -1999 -58 -1983 58
rect -2049 -70 -1983 -58
rect -1953 58 -1887 70
rect -1953 -58 -1937 58
rect -1903 -58 -1887 58
rect -1953 -70 -1887 -58
rect -1857 58 -1791 70
rect -1857 -58 -1841 58
rect -1807 -58 -1791 58
rect -1857 -70 -1791 -58
rect -1761 58 -1695 70
rect -1761 -58 -1745 58
rect -1711 -58 -1695 58
rect -1761 -70 -1695 -58
rect -1665 58 -1599 70
rect -1665 -58 -1649 58
rect -1615 -58 -1599 58
rect -1665 -70 -1599 -58
rect -1569 58 -1503 70
rect -1569 -58 -1553 58
rect -1519 -58 -1503 58
rect -1569 -70 -1503 -58
rect -1473 58 -1407 70
rect -1473 -58 -1457 58
rect -1423 -58 -1407 58
rect -1473 -70 -1407 -58
rect -1377 58 -1311 70
rect -1377 -58 -1361 58
rect -1327 -58 -1311 58
rect -1377 -70 -1311 -58
rect -1281 58 -1215 70
rect -1281 -58 -1265 58
rect -1231 -58 -1215 58
rect -1281 -70 -1215 -58
rect -1185 58 -1119 70
rect -1185 -58 -1169 58
rect -1135 -58 -1119 58
rect -1185 -70 -1119 -58
rect -1089 58 -1023 70
rect -1089 -58 -1073 58
rect -1039 -58 -1023 58
rect -1089 -70 -1023 -58
rect -993 58 -927 70
rect -993 -58 -977 58
rect -943 -58 -927 58
rect -993 -70 -927 -58
rect -897 58 -831 70
rect -897 -58 -881 58
rect -847 -58 -831 58
rect -897 -70 -831 -58
rect -801 58 -735 70
rect -801 -58 -785 58
rect -751 -58 -735 58
rect -801 -70 -735 -58
rect -705 58 -639 70
rect -705 -58 -689 58
rect -655 -58 -639 58
rect -705 -70 -639 -58
rect -609 58 -543 70
rect -609 -58 -593 58
rect -559 -58 -543 58
rect -609 -70 -543 -58
rect -513 58 -447 70
rect -513 -58 -497 58
rect -463 -58 -447 58
rect -513 -70 -447 -58
rect -417 58 -351 70
rect -417 -58 -401 58
rect -367 -58 -351 58
rect -417 -70 -351 -58
rect -321 58 -255 70
rect -321 -58 -305 58
rect -271 -58 -255 58
rect -321 -70 -255 -58
rect -225 58 -159 70
rect -225 -58 -209 58
rect -175 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 175 58
rect 209 -58 225 58
rect 159 -70 225 -58
rect 255 58 321 70
rect 255 -58 271 58
rect 305 -58 321 58
rect 255 -70 321 -58
rect 351 58 417 70
rect 351 -58 367 58
rect 401 -58 417 58
rect 351 -70 417 -58
rect 447 58 513 70
rect 447 -58 463 58
rect 497 -58 513 58
rect 447 -70 513 -58
rect 543 58 609 70
rect 543 -58 559 58
rect 593 -58 609 58
rect 543 -70 609 -58
rect 639 58 705 70
rect 639 -58 655 58
rect 689 -58 705 58
rect 639 -70 705 -58
rect 735 58 801 70
rect 735 -58 751 58
rect 785 -58 801 58
rect 735 -70 801 -58
rect 831 58 897 70
rect 831 -58 847 58
rect 881 -58 897 58
rect 831 -70 897 -58
rect 927 58 993 70
rect 927 -58 943 58
rect 977 -58 993 58
rect 927 -70 993 -58
rect 1023 58 1089 70
rect 1023 -58 1039 58
rect 1073 -58 1089 58
rect 1023 -70 1089 -58
rect 1119 58 1185 70
rect 1119 -58 1135 58
rect 1169 -58 1185 58
rect 1119 -70 1185 -58
rect 1215 58 1281 70
rect 1215 -58 1231 58
rect 1265 -58 1281 58
rect 1215 -70 1281 -58
rect 1311 58 1377 70
rect 1311 -58 1327 58
rect 1361 -58 1377 58
rect 1311 -70 1377 -58
rect 1407 58 1473 70
rect 1407 -58 1423 58
rect 1457 -58 1473 58
rect 1407 -70 1473 -58
rect 1503 58 1569 70
rect 1503 -58 1519 58
rect 1553 -58 1569 58
rect 1503 -70 1569 -58
rect 1599 58 1665 70
rect 1599 -58 1615 58
rect 1649 -58 1665 58
rect 1599 -70 1665 -58
rect 1695 58 1761 70
rect 1695 -58 1711 58
rect 1745 -58 1761 58
rect 1695 -70 1761 -58
rect 1791 58 1857 70
rect 1791 -58 1807 58
rect 1841 -58 1857 58
rect 1791 -70 1857 -58
rect 1887 58 1953 70
rect 1887 -58 1903 58
rect 1937 -58 1953 58
rect 1887 -70 1953 -58
rect 1983 58 2049 70
rect 1983 -58 1999 58
rect 2033 -58 2049 58
rect 1983 -70 2049 -58
rect 2079 58 2145 70
rect 2079 -58 2095 58
rect 2129 -58 2145 58
rect 2079 -70 2145 -58
rect 2175 58 2241 70
rect 2175 -58 2191 58
rect 2225 -58 2241 58
rect 2175 -70 2241 -58
rect 2271 58 2337 70
rect 2271 -58 2287 58
rect 2321 -58 2337 58
rect 2271 -70 2337 -58
rect 2367 58 2433 70
rect 2367 -58 2383 58
rect 2417 -58 2433 58
rect 2367 -70 2433 -58
rect 2463 58 2529 70
rect 2463 -58 2479 58
rect 2513 -58 2529 58
rect 2463 -70 2529 -58
rect 2559 58 2621 70
rect 2559 -58 2575 58
rect 2609 -58 2621 58
rect 2559 -70 2621 -58
<< pdiffc >>
rect -2609 -58 -2575 58
rect -2513 -58 -2479 58
rect -2417 -58 -2383 58
rect -2321 -58 -2287 58
rect -2225 -58 -2191 58
rect -2129 -58 -2095 58
rect -2033 -58 -1999 58
rect -1937 -58 -1903 58
rect -1841 -58 -1807 58
rect -1745 -58 -1711 58
rect -1649 -58 -1615 58
rect -1553 -58 -1519 58
rect -1457 -58 -1423 58
rect -1361 -58 -1327 58
rect -1265 -58 -1231 58
rect -1169 -58 -1135 58
rect -1073 -58 -1039 58
rect -977 -58 -943 58
rect -881 -58 -847 58
rect -785 -58 -751 58
rect -689 -58 -655 58
rect -593 -58 -559 58
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
rect 559 -58 593 58
rect 655 -58 689 58
rect 751 -58 785 58
rect 847 -58 881 58
rect 943 -58 977 58
rect 1039 -58 1073 58
rect 1135 -58 1169 58
rect 1231 -58 1265 58
rect 1327 -58 1361 58
rect 1423 -58 1457 58
rect 1519 -58 1553 58
rect 1615 -58 1649 58
rect 1711 -58 1745 58
rect 1807 -58 1841 58
rect 1903 -58 1937 58
rect 1999 -58 2033 58
rect 2095 -58 2129 58
rect 2191 -58 2225 58
rect 2287 -58 2321 58
rect 2383 -58 2417 58
rect 2479 -58 2513 58
rect 2575 -58 2609 58
<< nsubdiff >>
rect -2723 219 -2627 253
rect 2627 219 2723 253
rect -2723 157 -2689 219
rect 2689 157 2723 219
rect -2723 -219 -2689 -157
rect 2689 -219 2723 -157
rect -2723 -253 -2627 -219
rect 2627 -253 2723 -219
<< nsubdiffcont >>
rect -2627 219 2627 253
rect -2723 -157 -2689 157
rect 2689 -157 2723 157
rect -2627 -253 2627 -219
<< poly >>
rect -2481 151 -2415 167
rect -2481 117 -2465 151
rect -2431 117 -2415 151
rect -2481 101 -2415 117
rect -2289 151 -2223 167
rect -2289 117 -2273 151
rect -2239 117 -2223 151
rect -2289 101 -2223 117
rect -2097 151 -2031 167
rect -2097 117 -2081 151
rect -2047 117 -2031 151
rect -2097 101 -2031 117
rect -1905 151 -1839 167
rect -1905 117 -1889 151
rect -1855 117 -1839 151
rect -1905 101 -1839 117
rect -1713 151 -1647 167
rect -1713 117 -1697 151
rect -1663 117 -1647 151
rect -1713 101 -1647 117
rect -1521 151 -1455 167
rect -1521 117 -1505 151
rect -1471 117 -1455 151
rect -1521 101 -1455 117
rect -1329 151 -1263 167
rect -1329 117 -1313 151
rect -1279 117 -1263 151
rect -1329 101 -1263 117
rect -1137 151 -1071 167
rect -1137 117 -1121 151
rect -1087 117 -1071 151
rect -1137 101 -1071 117
rect -945 151 -879 167
rect -945 117 -929 151
rect -895 117 -879 151
rect -945 101 -879 117
rect -753 151 -687 167
rect -753 117 -737 151
rect -703 117 -687 151
rect -753 101 -687 117
rect -561 151 -495 167
rect -561 117 -545 151
rect -511 117 -495 151
rect -561 101 -495 117
rect -369 151 -303 167
rect -369 117 -353 151
rect -319 117 -303 151
rect -369 101 -303 117
rect -177 151 -111 167
rect -177 117 -161 151
rect -127 117 -111 151
rect -177 101 -111 117
rect 15 151 81 167
rect 15 117 31 151
rect 65 117 81 151
rect 15 101 81 117
rect 207 151 273 167
rect 207 117 223 151
rect 257 117 273 151
rect 207 101 273 117
rect 399 151 465 167
rect 399 117 415 151
rect 449 117 465 151
rect 399 101 465 117
rect 591 151 657 167
rect 591 117 607 151
rect 641 117 657 151
rect 591 101 657 117
rect 783 151 849 167
rect 783 117 799 151
rect 833 117 849 151
rect 783 101 849 117
rect 975 151 1041 167
rect 975 117 991 151
rect 1025 117 1041 151
rect 975 101 1041 117
rect 1167 151 1233 167
rect 1167 117 1183 151
rect 1217 117 1233 151
rect 1167 101 1233 117
rect 1359 151 1425 167
rect 1359 117 1375 151
rect 1409 117 1425 151
rect 1359 101 1425 117
rect 1551 151 1617 167
rect 1551 117 1567 151
rect 1601 117 1617 151
rect 1551 101 1617 117
rect 1743 151 1809 167
rect 1743 117 1759 151
rect 1793 117 1809 151
rect 1743 101 1809 117
rect 1935 151 2001 167
rect 1935 117 1951 151
rect 1985 117 2001 151
rect 1935 101 2001 117
rect 2127 151 2193 167
rect 2127 117 2143 151
rect 2177 117 2193 151
rect 2127 101 2193 117
rect 2319 151 2385 167
rect 2319 117 2335 151
rect 2369 117 2385 151
rect 2319 101 2385 117
rect 2511 151 2577 167
rect 2511 117 2527 151
rect 2561 117 2577 151
rect 2511 101 2577 117
rect -2559 70 -2529 96
rect -2463 70 -2433 101
rect -2367 70 -2337 96
rect -2271 70 -2241 101
rect -2175 70 -2145 96
rect -2079 70 -2049 101
rect -1983 70 -1953 96
rect -1887 70 -1857 101
rect -1791 70 -1761 96
rect -1695 70 -1665 101
rect -1599 70 -1569 96
rect -1503 70 -1473 101
rect -1407 70 -1377 96
rect -1311 70 -1281 101
rect -1215 70 -1185 96
rect -1119 70 -1089 101
rect -1023 70 -993 96
rect -927 70 -897 101
rect -831 70 -801 96
rect -735 70 -705 101
rect -639 70 -609 96
rect -543 70 -513 101
rect -447 70 -417 96
rect -351 70 -321 101
rect -255 70 -225 96
rect -159 70 -129 101
rect -63 70 -33 96
rect 33 70 63 101
rect 129 70 159 96
rect 225 70 255 101
rect 321 70 351 96
rect 417 70 447 101
rect 513 70 543 96
rect 609 70 639 101
rect 705 70 735 96
rect 801 70 831 101
rect 897 70 927 96
rect 993 70 1023 101
rect 1089 70 1119 96
rect 1185 70 1215 101
rect 1281 70 1311 96
rect 1377 70 1407 101
rect 1473 70 1503 96
rect 1569 70 1599 101
rect 1665 70 1695 96
rect 1761 70 1791 101
rect 1857 70 1887 96
rect 1953 70 1983 101
rect 2049 70 2079 96
rect 2145 70 2175 101
rect 2241 70 2271 96
rect 2337 70 2367 101
rect 2433 70 2463 96
rect 2529 70 2559 101
rect -2559 -101 -2529 -70
rect -2463 -96 -2433 -70
rect -2367 -101 -2337 -70
rect -2271 -96 -2241 -70
rect -2175 -101 -2145 -70
rect -2079 -96 -2049 -70
rect -1983 -101 -1953 -70
rect -1887 -96 -1857 -70
rect -1791 -101 -1761 -70
rect -1695 -96 -1665 -70
rect -1599 -101 -1569 -70
rect -1503 -96 -1473 -70
rect -1407 -101 -1377 -70
rect -1311 -96 -1281 -70
rect -1215 -101 -1185 -70
rect -1119 -96 -1089 -70
rect -1023 -101 -993 -70
rect -927 -96 -897 -70
rect -831 -101 -801 -70
rect -735 -96 -705 -70
rect -639 -101 -609 -70
rect -543 -96 -513 -70
rect -447 -101 -417 -70
rect -351 -96 -321 -70
rect -255 -101 -225 -70
rect -159 -96 -129 -70
rect -63 -101 -33 -70
rect 33 -96 63 -70
rect 129 -101 159 -70
rect 225 -96 255 -70
rect 321 -101 351 -70
rect 417 -96 447 -70
rect 513 -101 543 -70
rect 609 -96 639 -70
rect 705 -101 735 -70
rect 801 -96 831 -70
rect 897 -101 927 -70
rect 993 -96 1023 -70
rect 1089 -101 1119 -70
rect 1185 -96 1215 -70
rect 1281 -101 1311 -70
rect 1377 -96 1407 -70
rect 1473 -101 1503 -70
rect 1569 -96 1599 -70
rect 1665 -101 1695 -70
rect 1761 -96 1791 -70
rect 1857 -101 1887 -70
rect 1953 -96 1983 -70
rect 2049 -101 2079 -70
rect 2145 -96 2175 -70
rect 2241 -101 2271 -70
rect 2337 -96 2367 -70
rect 2433 -101 2463 -70
rect 2529 -96 2559 -70
rect -2577 -117 -2511 -101
rect -2577 -151 -2561 -117
rect -2527 -151 -2511 -117
rect -2577 -167 -2511 -151
rect -2385 -117 -2319 -101
rect -2385 -151 -2369 -117
rect -2335 -151 -2319 -117
rect -2385 -167 -2319 -151
rect -2193 -117 -2127 -101
rect -2193 -151 -2177 -117
rect -2143 -151 -2127 -117
rect -2193 -167 -2127 -151
rect -2001 -117 -1935 -101
rect -2001 -151 -1985 -117
rect -1951 -151 -1935 -117
rect -2001 -167 -1935 -151
rect -1809 -117 -1743 -101
rect -1809 -151 -1793 -117
rect -1759 -151 -1743 -117
rect -1809 -167 -1743 -151
rect -1617 -117 -1551 -101
rect -1617 -151 -1601 -117
rect -1567 -151 -1551 -117
rect -1617 -167 -1551 -151
rect -1425 -117 -1359 -101
rect -1425 -151 -1409 -117
rect -1375 -151 -1359 -117
rect -1425 -167 -1359 -151
rect -1233 -117 -1167 -101
rect -1233 -151 -1217 -117
rect -1183 -151 -1167 -117
rect -1233 -167 -1167 -151
rect -1041 -117 -975 -101
rect -1041 -151 -1025 -117
rect -991 -151 -975 -117
rect -1041 -167 -975 -151
rect -849 -117 -783 -101
rect -849 -151 -833 -117
rect -799 -151 -783 -117
rect -849 -167 -783 -151
rect -657 -117 -591 -101
rect -657 -151 -641 -117
rect -607 -151 -591 -117
rect -657 -167 -591 -151
rect -465 -117 -399 -101
rect -465 -151 -449 -117
rect -415 -151 -399 -117
rect -465 -167 -399 -151
rect -273 -117 -207 -101
rect -273 -151 -257 -117
rect -223 -151 -207 -117
rect -273 -167 -207 -151
rect -81 -117 -15 -101
rect -81 -151 -65 -117
rect -31 -151 -15 -117
rect -81 -167 -15 -151
rect 111 -117 177 -101
rect 111 -151 127 -117
rect 161 -151 177 -117
rect 111 -167 177 -151
rect 303 -117 369 -101
rect 303 -151 319 -117
rect 353 -151 369 -117
rect 303 -167 369 -151
rect 495 -117 561 -101
rect 495 -151 511 -117
rect 545 -151 561 -117
rect 495 -167 561 -151
rect 687 -117 753 -101
rect 687 -151 703 -117
rect 737 -151 753 -117
rect 687 -167 753 -151
rect 879 -117 945 -101
rect 879 -151 895 -117
rect 929 -151 945 -117
rect 879 -167 945 -151
rect 1071 -117 1137 -101
rect 1071 -151 1087 -117
rect 1121 -151 1137 -117
rect 1071 -167 1137 -151
rect 1263 -117 1329 -101
rect 1263 -151 1279 -117
rect 1313 -151 1329 -117
rect 1263 -167 1329 -151
rect 1455 -117 1521 -101
rect 1455 -151 1471 -117
rect 1505 -151 1521 -117
rect 1455 -167 1521 -151
rect 1647 -117 1713 -101
rect 1647 -151 1663 -117
rect 1697 -151 1713 -117
rect 1647 -167 1713 -151
rect 1839 -117 1905 -101
rect 1839 -151 1855 -117
rect 1889 -151 1905 -117
rect 1839 -167 1905 -151
rect 2031 -117 2097 -101
rect 2031 -151 2047 -117
rect 2081 -151 2097 -117
rect 2031 -167 2097 -151
rect 2223 -117 2289 -101
rect 2223 -151 2239 -117
rect 2273 -151 2289 -117
rect 2223 -167 2289 -151
rect 2415 -117 2481 -101
rect 2415 -151 2431 -117
rect 2465 -151 2481 -117
rect 2415 -167 2481 -151
<< polycont >>
rect -2465 117 -2431 151
rect -2273 117 -2239 151
rect -2081 117 -2047 151
rect -1889 117 -1855 151
rect -1697 117 -1663 151
rect -1505 117 -1471 151
rect -1313 117 -1279 151
rect -1121 117 -1087 151
rect -929 117 -895 151
rect -737 117 -703 151
rect -545 117 -511 151
rect -353 117 -319 151
rect -161 117 -127 151
rect 31 117 65 151
rect 223 117 257 151
rect 415 117 449 151
rect 607 117 641 151
rect 799 117 833 151
rect 991 117 1025 151
rect 1183 117 1217 151
rect 1375 117 1409 151
rect 1567 117 1601 151
rect 1759 117 1793 151
rect 1951 117 1985 151
rect 2143 117 2177 151
rect 2335 117 2369 151
rect 2527 117 2561 151
rect -2561 -151 -2527 -117
rect -2369 -151 -2335 -117
rect -2177 -151 -2143 -117
rect -1985 -151 -1951 -117
rect -1793 -151 -1759 -117
rect -1601 -151 -1567 -117
rect -1409 -151 -1375 -117
rect -1217 -151 -1183 -117
rect -1025 -151 -991 -117
rect -833 -151 -799 -117
rect -641 -151 -607 -117
rect -449 -151 -415 -117
rect -257 -151 -223 -117
rect -65 -151 -31 -117
rect 127 -151 161 -117
rect 319 -151 353 -117
rect 511 -151 545 -117
rect 703 -151 737 -117
rect 895 -151 929 -117
rect 1087 -151 1121 -117
rect 1279 -151 1313 -117
rect 1471 -151 1505 -117
rect 1663 -151 1697 -117
rect 1855 -151 1889 -117
rect 2047 -151 2081 -117
rect 2239 -151 2273 -117
rect 2431 -151 2465 -117
<< locali >>
rect -2723 219 -2627 253
rect 2627 219 2723 253
rect -2723 157 -2689 219
rect 2689 157 2723 219
rect -2481 117 -2465 151
rect -2431 117 -2415 151
rect -2289 117 -2273 151
rect -2239 117 -2223 151
rect -2097 117 -2081 151
rect -2047 117 -2031 151
rect -1905 117 -1889 151
rect -1855 117 -1839 151
rect -1713 117 -1697 151
rect -1663 117 -1647 151
rect -1521 117 -1505 151
rect -1471 117 -1455 151
rect -1329 117 -1313 151
rect -1279 117 -1263 151
rect -1137 117 -1121 151
rect -1087 117 -1071 151
rect -945 117 -929 151
rect -895 117 -879 151
rect -753 117 -737 151
rect -703 117 -687 151
rect -561 117 -545 151
rect -511 117 -495 151
rect -369 117 -353 151
rect -319 117 -303 151
rect -177 117 -161 151
rect -127 117 -111 151
rect 15 117 31 151
rect 65 117 81 151
rect 207 117 223 151
rect 257 117 273 151
rect 399 117 415 151
rect 449 117 465 151
rect 591 117 607 151
rect 641 117 657 151
rect 783 117 799 151
rect 833 117 849 151
rect 975 117 991 151
rect 1025 117 1041 151
rect 1167 117 1183 151
rect 1217 117 1233 151
rect 1359 117 1375 151
rect 1409 117 1425 151
rect 1551 117 1567 151
rect 1601 117 1617 151
rect 1743 117 1759 151
rect 1793 117 1809 151
rect 1935 117 1951 151
rect 1985 117 2001 151
rect 2127 117 2143 151
rect 2177 117 2193 151
rect 2319 117 2335 151
rect 2369 117 2385 151
rect 2511 117 2527 151
rect 2561 117 2577 151
rect -2609 58 -2575 74
rect -2609 -74 -2575 -58
rect -2513 58 -2479 74
rect -2513 -74 -2479 -58
rect -2417 58 -2383 74
rect -2417 -74 -2383 -58
rect -2321 58 -2287 74
rect -2321 -74 -2287 -58
rect -2225 58 -2191 74
rect -2225 -74 -2191 -58
rect -2129 58 -2095 74
rect -2129 -74 -2095 -58
rect -2033 58 -1999 74
rect -2033 -74 -1999 -58
rect -1937 58 -1903 74
rect -1937 -74 -1903 -58
rect -1841 58 -1807 74
rect -1841 -74 -1807 -58
rect -1745 58 -1711 74
rect -1745 -74 -1711 -58
rect -1649 58 -1615 74
rect -1649 -74 -1615 -58
rect -1553 58 -1519 74
rect -1553 -74 -1519 -58
rect -1457 58 -1423 74
rect -1457 -74 -1423 -58
rect -1361 58 -1327 74
rect -1361 -74 -1327 -58
rect -1265 58 -1231 74
rect -1265 -74 -1231 -58
rect -1169 58 -1135 74
rect -1169 -74 -1135 -58
rect -1073 58 -1039 74
rect -1073 -74 -1039 -58
rect -977 58 -943 74
rect -977 -74 -943 -58
rect -881 58 -847 74
rect -881 -74 -847 -58
rect -785 58 -751 74
rect -785 -74 -751 -58
rect -689 58 -655 74
rect -689 -74 -655 -58
rect -593 58 -559 74
rect -593 -74 -559 -58
rect -497 58 -463 74
rect -497 -74 -463 -58
rect -401 58 -367 74
rect -401 -74 -367 -58
rect -305 58 -271 74
rect -305 -74 -271 -58
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect 271 58 305 74
rect 271 -74 305 -58
rect 367 58 401 74
rect 367 -74 401 -58
rect 463 58 497 74
rect 463 -74 497 -58
rect 559 58 593 74
rect 559 -74 593 -58
rect 655 58 689 74
rect 655 -74 689 -58
rect 751 58 785 74
rect 751 -74 785 -58
rect 847 58 881 74
rect 847 -74 881 -58
rect 943 58 977 74
rect 943 -74 977 -58
rect 1039 58 1073 74
rect 1039 -74 1073 -58
rect 1135 58 1169 74
rect 1135 -74 1169 -58
rect 1231 58 1265 74
rect 1231 -74 1265 -58
rect 1327 58 1361 74
rect 1327 -74 1361 -58
rect 1423 58 1457 74
rect 1423 -74 1457 -58
rect 1519 58 1553 74
rect 1519 -74 1553 -58
rect 1615 58 1649 74
rect 1615 -74 1649 -58
rect 1711 58 1745 74
rect 1711 -74 1745 -58
rect 1807 58 1841 74
rect 1807 -74 1841 -58
rect 1903 58 1937 74
rect 1903 -74 1937 -58
rect 1999 58 2033 74
rect 1999 -74 2033 -58
rect 2095 58 2129 74
rect 2095 -74 2129 -58
rect 2191 58 2225 74
rect 2191 -74 2225 -58
rect 2287 58 2321 74
rect 2287 -74 2321 -58
rect 2383 58 2417 74
rect 2383 -74 2417 -58
rect 2479 58 2513 74
rect 2479 -74 2513 -58
rect 2575 58 2609 74
rect 2575 -74 2609 -58
rect -2577 -151 -2561 -117
rect -2527 -151 -2511 -117
rect -2385 -151 -2369 -117
rect -2335 -151 -2319 -117
rect -2193 -151 -2177 -117
rect -2143 -151 -2127 -117
rect -2001 -151 -1985 -117
rect -1951 -151 -1935 -117
rect -1809 -151 -1793 -117
rect -1759 -151 -1743 -117
rect -1617 -151 -1601 -117
rect -1567 -151 -1551 -117
rect -1425 -151 -1409 -117
rect -1375 -151 -1359 -117
rect -1233 -151 -1217 -117
rect -1183 -151 -1167 -117
rect -1041 -151 -1025 -117
rect -991 -151 -975 -117
rect -849 -151 -833 -117
rect -799 -151 -783 -117
rect -657 -151 -641 -117
rect -607 -151 -591 -117
rect -465 -151 -449 -117
rect -415 -151 -399 -117
rect -273 -151 -257 -117
rect -223 -151 -207 -117
rect -81 -151 -65 -117
rect -31 -151 -15 -117
rect 111 -151 127 -117
rect 161 -151 177 -117
rect 303 -151 319 -117
rect 353 -151 369 -117
rect 495 -151 511 -117
rect 545 -151 561 -117
rect 687 -151 703 -117
rect 737 -151 753 -117
rect 879 -151 895 -117
rect 929 -151 945 -117
rect 1071 -151 1087 -117
rect 1121 -151 1137 -117
rect 1263 -151 1279 -117
rect 1313 -151 1329 -117
rect 1455 -151 1471 -117
rect 1505 -151 1521 -117
rect 1647 -151 1663 -117
rect 1697 -151 1713 -117
rect 1839 -151 1855 -117
rect 1889 -151 1905 -117
rect 2031 -151 2047 -117
rect 2081 -151 2097 -117
rect 2223 -151 2239 -117
rect 2273 -151 2289 -117
rect 2415 -151 2431 -117
rect 2465 -151 2481 -117
rect -2723 -219 -2689 -157
rect 2689 -219 2723 -157
rect -2723 -253 -2627 -219
rect 2627 -253 2723 -219
<< viali >>
rect -2465 117 -2431 151
rect -2273 117 -2239 151
rect -2081 117 -2047 151
rect -1889 117 -1855 151
rect -1697 117 -1663 151
rect -1505 117 -1471 151
rect -1313 117 -1279 151
rect -1121 117 -1087 151
rect -929 117 -895 151
rect -737 117 -703 151
rect -545 117 -511 151
rect -353 117 -319 151
rect -161 117 -127 151
rect 31 117 65 151
rect 223 117 257 151
rect 415 117 449 151
rect 607 117 641 151
rect 799 117 833 151
rect 991 117 1025 151
rect 1183 117 1217 151
rect 1375 117 1409 151
rect 1567 117 1601 151
rect 1759 117 1793 151
rect 1951 117 1985 151
rect 2143 117 2177 151
rect 2335 117 2369 151
rect 2527 117 2561 151
rect -2609 -58 -2575 58
rect -2513 -58 -2479 58
rect -2417 -58 -2383 58
rect -2321 -58 -2287 58
rect -2225 -58 -2191 58
rect -2129 -58 -2095 58
rect -2033 -58 -1999 58
rect -1937 -58 -1903 58
rect -1841 -58 -1807 58
rect -1745 -58 -1711 58
rect -1649 -58 -1615 58
rect -1553 -58 -1519 58
rect -1457 -58 -1423 58
rect -1361 -58 -1327 58
rect -1265 -58 -1231 58
rect -1169 -58 -1135 58
rect -1073 -58 -1039 58
rect -977 -58 -943 58
rect -881 -58 -847 58
rect -785 -58 -751 58
rect -689 -58 -655 58
rect -593 -58 -559 58
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
rect 559 -58 593 58
rect 655 -58 689 58
rect 751 -58 785 58
rect 847 -58 881 58
rect 943 -58 977 58
rect 1039 -58 1073 58
rect 1135 -58 1169 58
rect 1231 -58 1265 58
rect 1327 -58 1361 58
rect 1423 -58 1457 58
rect 1519 -58 1553 58
rect 1615 -58 1649 58
rect 1711 -58 1745 58
rect 1807 -58 1841 58
rect 1903 -58 1937 58
rect 1999 -58 2033 58
rect 2095 -58 2129 58
rect 2191 -58 2225 58
rect 2287 -58 2321 58
rect 2383 -58 2417 58
rect 2479 -58 2513 58
rect 2575 -58 2609 58
rect -2561 -151 -2527 -117
rect -2369 -151 -2335 -117
rect -2177 -151 -2143 -117
rect -1985 -151 -1951 -117
rect -1793 -151 -1759 -117
rect -1601 -151 -1567 -117
rect -1409 -151 -1375 -117
rect -1217 -151 -1183 -117
rect -1025 -151 -991 -117
rect -833 -151 -799 -117
rect -641 -151 -607 -117
rect -449 -151 -415 -117
rect -257 -151 -223 -117
rect -65 -151 -31 -117
rect 127 -151 161 -117
rect 319 -151 353 -117
rect 511 -151 545 -117
rect 703 -151 737 -117
rect 895 -151 929 -117
rect 1087 -151 1121 -117
rect 1279 -151 1313 -117
rect 1471 -151 1505 -117
rect 1663 -151 1697 -117
rect 1855 -151 1889 -117
rect 2047 -151 2081 -117
rect 2239 -151 2273 -117
rect 2431 -151 2465 -117
<< metal1 >>
rect -2477 151 -2419 157
rect -2477 117 -2465 151
rect -2431 117 -2419 151
rect -2477 111 -2419 117
rect -2285 151 -2227 157
rect -2285 117 -2273 151
rect -2239 117 -2227 151
rect -2285 111 -2227 117
rect -2093 151 -2035 157
rect -2093 117 -2081 151
rect -2047 117 -2035 151
rect -2093 111 -2035 117
rect -1901 151 -1843 157
rect -1901 117 -1889 151
rect -1855 117 -1843 151
rect -1901 111 -1843 117
rect -1709 151 -1651 157
rect -1709 117 -1697 151
rect -1663 117 -1651 151
rect -1709 111 -1651 117
rect -1517 151 -1459 157
rect -1517 117 -1505 151
rect -1471 117 -1459 151
rect -1517 111 -1459 117
rect -1325 151 -1267 157
rect -1325 117 -1313 151
rect -1279 117 -1267 151
rect -1325 111 -1267 117
rect -1133 151 -1075 157
rect -1133 117 -1121 151
rect -1087 117 -1075 151
rect -1133 111 -1075 117
rect -941 151 -883 157
rect -941 117 -929 151
rect -895 117 -883 151
rect -941 111 -883 117
rect -749 151 -691 157
rect -749 117 -737 151
rect -703 117 -691 151
rect -749 111 -691 117
rect -557 151 -499 157
rect -557 117 -545 151
rect -511 117 -499 151
rect -557 111 -499 117
rect -365 151 -307 157
rect -365 117 -353 151
rect -319 117 -307 151
rect -365 111 -307 117
rect -173 151 -115 157
rect -173 117 -161 151
rect -127 117 -115 151
rect -173 111 -115 117
rect 19 151 77 157
rect 19 117 31 151
rect 65 117 77 151
rect 19 111 77 117
rect 211 151 269 157
rect 211 117 223 151
rect 257 117 269 151
rect 211 111 269 117
rect 403 151 461 157
rect 403 117 415 151
rect 449 117 461 151
rect 403 111 461 117
rect 595 151 653 157
rect 595 117 607 151
rect 641 117 653 151
rect 595 111 653 117
rect 787 151 845 157
rect 787 117 799 151
rect 833 117 845 151
rect 787 111 845 117
rect 979 151 1037 157
rect 979 117 991 151
rect 1025 117 1037 151
rect 979 111 1037 117
rect 1171 151 1229 157
rect 1171 117 1183 151
rect 1217 117 1229 151
rect 1171 111 1229 117
rect 1363 151 1421 157
rect 1363 117 1375 151
rect 1409 117 1421 151
rect 1363 111 1421 117
rect 1555 151 1613 157
rect 1555 117 1567 151
rect 1601 117 1613 151
rect 1555 111 1613 117
rect 1747 151 1805 157
rect 1747 117 1759 151
rect 1793 117 1805 151
rect 1747 111 1805 117
rect 1939 151 1997 157
rect 1939 117 1951 151
rect 1985 117 1997 151
rect 1939 111 1997 117
rect 2131 151 2189 157
rect 2131 117 2143 151
rect 2177 117 2189 151
rect 2131 111 2189 117
rect 2323 151 2381 157
rect 2323 117 2335 151
rect 2369 117 2381 151
rect 2323 111 2381 117
rect 2515 151 2573 157
rect 2515 117 2527 151
rect 2561 117 2573 151
rect 2515 111 2573 117
rect -2615 58 -2569 70
rect -2615 -58 -2609 58
rect -2575 -58 -2569 58
rect -2615 -70 -2569 -58
rect -2519 58 -2473 70
rect -2519 -58 -2513 58
rect -2479 -58 -2473 58
rect -2519 -70 -2473 -58
rect -2423 58 -2377 70
rect -2423 -58 -2417 58
rect -2383 -58 -2377 58
rect -2423 -70 -2377 -58
rect -2327 58 -2281 70
rect -2327 -58 -2321 58
rect -2287 -58 -2281 58
rect -2327 -70 -2281 -58
rect -2231 58 -2185 70
rect -2231 -58 -2225 58
rect -2191 -58 -2185 58
rect -2231 -70 -2185 -58
rect -2135 58 -2089 70
rect -2135 -58 -2129 58
rect -2095 -58 -2089 58
rect -2135 -70 -2089 -58
rect -2039 58 -1993 70
rect -2039 -58 -2033 58
rect -1999 -58 -1993 58
rect -2039 -70 -1993 -58
rect -1943 58 -1897 70
rect -1943 -58 -1937 58
rect -1903 -58 -1897 58
rect -1943 -70 -1897 -58
rect -1847 58 -1801 70
rect -1847 -58 -1841 58
rect -1807 -58 -1801 58
rect -1847 -70 -1801 -58
rect -1751 58 -1705 70
rect -1751 -58 -1745 58
rect -1711 -58 -1705 58
rect -1751 -70 -1705 -58
rect -1655 58 -1609 70
rect -1655 -58 -1649 58
rect -1615 -58 -1609 58
rect -1655 -70 -1609 -58
rect -1559 58 -1513 70
rect -1559 -58 -1553 58
rect -1519 -58 -1513 58
rect -1559 -70 -1513 -58
rect -1463 58 -1417 70
rect -1463 -58 -1457 58
rect -1423 -58 -1417 58
rect -1463 -70 -1417 -58
rect -1367 58 -1321 70
rect -1367 -58 -1361 58
rect -1327 -58 -1321 58
rect -1367 -70 -1321 -58
rect -1271 58 -1225 70
rect -1271 -58 -1265 58
rect -1231 -58 -1225 58
rect -1271 -70 -1225 -58
rect -1175 58 -1129 70
rect -1175 -58 -1169 58
rect -1135 -58 -1129 58
rect -1175 -70 -1129 -58
rect -1079 58 -1033 70
rect -1079 -58 -1073 58
rect -1039 -58 -1033 58
rect -1079 -70 -1033 -58
rect -983 58 -937 70
rect -983 -58 -977 58
rect -943 -58 -937 58
rect -983 -70 -937 -58
rect -887 58 -841 70
rect -887 -58 -881 58
rect -847 -58 -841 58
rect -887 -70 -841 -58
rect -791 58 -745 70
rect -791 -58 -785 58
rect -751 -58 -745 58
rect -791 -70 -745 -58
rect -695 58 -649 70
rect -695 -58 -689 58
rect -655 -58 -649 58
rect -695 -70 -649 -58
rect -599 58 -553 70
rect -599 -58 -593 58
rect -559 -58 -553 58
rect -599 -70 -553 -58
rect -503 58 -457 70
rect -503 -58 -497 58
rect -463 -58 -457 58
rect -503 -70 -457 -58
rect -407 58 -361 70
rect -407 -58 -401 58
rect -367 -58 -361 58
rect -407 -70 -361 -58
rect -311 58 -265 70
rect -311 -58 -305 58
rect -271 -58 -265 58
rect -311 -70 -265 -58
rect -215 58 -169 70
rect -215 -58 -209 58
rect -175 -58 -169 58
rect -215 -70 -169 -58
rect -119 58 -73 70
rect -119 -58 -113 58
rect -79 -58 -73 58
rect -119 -70 -73 -58
rect -23 58 23 70
rect -23 -58 -17 58
rect 17 -58 23 58
rect -23 -70 23 -58
rect 73 58 119 70
rect 73 -58 79 58
rect 113 -58 119 58
rect 73 -70 119 -58
rect 169 58 215 70
rect 169 -58 175 58
rect 209 -58 215 58
rect 169 -70 215 -58
rect 265 58 311 70
rect 265 -58 271 58
rect 305 -58 311 58
rect 265 -70 311 -58
rect 361 58 407 70
rect 361 -58 367 58
rect 401 -58 407 58
rect 361 -70 407 -58
rect 457 58 503 70
rect 457 -58 463 58
rect 497 -58 503 58
rect 457 -70 503 -58
rect 553 58 599 70
rect 553 -58 559 58
rect 593 -58 599 58
rect 553 -70 599 -58
rect 649 58 695 70
rect 649 -58 655 58
rect 689 -58 695 58
rect 649 -70 695 -58
rect 745 58 791 70
rect 745 -58 751 58
rect 785 -58 791 58
rect 745 -70 791 -58
rect 841 58 887 70
rect 841 -58 847 58
rect 881 -58 887 58
rect 841 -70 887 -58
rect 937 58 983 70
rect 937 -58 943 58
rect 977 -58 983 58
rect 937 -70 983 -58
rect 1033 58 1079 70
rect 1033 -58 1039 58
rect 1073 -58 1079 58
rect 1033 -70 1079 -58
rect 1129 58 1175 70
rect 1129 -58 1135 58
rect 1169 -58 1175 58
rect 1129 -70 1175 -58
rect 1225 58 1271 70
rect 1225 -58 1231 58
rect 1265 -58 1271 58
rect 1225 -70 1271 -58
rect 1321 58 1367 70
rect 1321 -58 1327 58
rect 1361 -58 1367 58
rect 1321 -70 1367 -58
rect 1417 58 1463 70
rect 1417 -58 1423 58
rect 1457 -58 1463 58
rect 1417 -70 1463 -58
rect 1513 58 1559 70
rect 1513 -58 1519 58
rect 1553 -58 1559 58
rect 1513 -70 1559 -58
rect 1609 58 1655 70
rect 1609 -58 1615 58
rect 1649 -58 1655 58
rect 1609 -70 1655 -58
rect 1705 58 1751 70
rect 1705 -58 1711 58
rect 1745 -58 1751 58
rect 1705 -70 1751 -58
rect 1801 58 1847 70
rect 1801 -58 1807 58
rect 1841 -58 1847 58
rect 1801 -70 1847 -58
rect 1897 58 1943 70
rect 1897 -58 1903 58
rect 1937 -58 1943 58
rect 1897 -70 1943 -58
rect 1993 58 2039 70
rect 1993 -58 1999 58
rect 2033 -58 2039 58
rect 1993 -70 2039 -58
rect 2089 58 2135 70
rect 2089 -58 2095 58
rect 2129 -58 2135 58
rect 2089 -70 2135 -58
rect 2185 58 2231 70
rect 2185 -58 2191 58
rect 2225 -58 2231 58
rect 2185 -70 2231 -58
rect 2281 58 2327 70
rect 2281 -58 2287 58
rect 2321 -58 2327 58
rect 2281 -70 2327 -58
rect 2377 58 2423 70
rect 2377 -58 2383 58
rect 2417 -58 2423 58
rect 2377 -70 2423 -58
rect 2473 58 2519 70
rect 2473 -58 2479 58
rect 2513 -58 2519 58
rect 2473 -70 2519 -58
rect 2569 58 2615 70
rect 2569 -58 2575 58
rect 2609 -58 2615 58
rect 2569 -70 2615 -58
rect -2573 -117 -2515 -111
rect -2573 -151 -2561 -117
rect -2527 -151 -2515 -117
rect -2573 -157 -2515 -151
rect -2381 -117 -2323 -111
rect -2381 -151 -2369 -117
rect -2335 -151 -2323 -117
rect -2381 -157 -2323 -151
rect -2189 -117 -2131 -111
rect -2189 -151 -2177 -117
rect -2143 -151 -2131 -117
rect -2189 -157 -2131 -151
rect -1997 -117 -1939 -111
rect -1997 -151 -1985 -117
rect -1951 -151 -1939 -117
rect -1997 -157 -1939 -151
rect -1805 -117 -1747 -111
rect -1805 -151 -1793 -117
rect -1759 -151 -1747 -117
rect -1805 -157 -1747 -151
rect -1613 -117 -1555 -111
rect -1613 -151 -1601 -117
rect -1567 -151 -1555 -117
rect -1613 -157 -1555 -151
rect -1421 -117 -1363 -111
rect -1421 -151 -1409 -117
rect -1375 -151 -1363 -117
rect -1421 -157 -1363 -151
rect -1229 -117 -1171 -111
rect -1229 -151 -1217 -117
rect -1183 -151 -1171 -117
rect -1229 -157 -1171 -151
rect -1037 -117 -979 -111
rect -1037 -151 -1025 -117
rect -991 -151 -979 -117
rect -1037 -157 -979 -151
rect -845 -117 -787 -111
rect -845 -151 -833 -117
rect -799 -151 -787 -117
rect -845 -157 -787 -151
rect -653 -117 -595 -111
rect -653 -151 -641 -117
rect -607 -151 -595 -117
rect -653 -157 -595 -151
rect -461 -117 -403 -111
rect -461 -151 -449 -117
rect -415 -151 -403 -117
rect -461 -157 -403 -151
rect -269 -117 -211 -111
rect -269 -151 -257 -117
rect -223 -151 -211 -117
rect -269 -157 -211 -151
rect -77 -117 -19 -111
rect -77 -151 -65 -117
rect -31 -151 -19 -117
rect -77 -157 -19 -151
rect 115 -117 173 -111
rect 115 -151 127 -117
rect 161 -151 173 -117
rect 115 -157 173 -151
rect 307 -117 365 -111
rect 307 -151 319 -117
rect 353 -151 365 -117
rect 307 -157 365 -151
rect 499 -117 557 -111
rect 499 -151 511 -117
rect 545 -151 557 -117
rect 499 -157 557 -151
rect 691 -117 749 -111
rect 691 -151 703 -117
rect 737 -151 749 -117
rect 691 -157 749 -151
rect 883 -117 941 -111
rect 883 -151 895 -117
rect 929 -151 941 -117
rect 883 -157 941 -151
rect 1075 -117 1133 -111
rect 1075 -151 1087 -117
rect 1121 -151 1133 -117
rect 1075 -157 1133 -151
rect 1267 -117 1325 -111
rect 1267 -151 1279 -117
rect 1313 -151 1325 -117
rect 1267 -157 1325 -151
rect 1459 -117 1517 -111
rect 1459 -151 1471 -117
rect 1505 -151 1517 -117
rect 1459 -157 1517 -151
rect 1651 -117 1709 -111
rect 1651 -151 1663 -117
rect 1697 -151 1709 -117
rect 1651 -157 1709 -151
rect 1843 -117 1901 -111
rect 1843 -151 1855 -117
rect 1889 -151 1901 -117
rect 1843 -157 1901 -151
rect 2035 -117 2093 -111
rect 2035 -151 2047 -117
rect 2081 -151 2093 -117
rect 2035 -157 2093 -151
rect 2227 -117 2285 -111
rect 2227 -151 2239 -117
rect 2273 -151 2285 -117
rect 2227 -157 2285 -151
rect 2419 -117 2477 -111
rect 2419 -151 2431 -117
rect 2465 -151 2477 -117
rect 2419 -157 2477 -151
<< properties >>
string FIXED_BBOX -2706 -236 2706 236
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.7 l 0.15 m 1 nf 54 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
