magic
tech sky130A
magscale 1 2
timestamp 1718283729
<< pwell >>
rect -201 -1482 201 1482
<< psubdiff >>
rect -165 1412 -69 1446
rect 69 1412 165 1446
rect -165 1350 -131 1412
rect 131 1350 165 1412
rect -165 -1412 -131 -1350
rect 131 -1412 165 -1350
rect -165 -1446 -69 -1412
rect 69 -1446 165 -1412
<< psubdiffcont >>
rect -69 1412 69 1446
rect -165 -1350 -131 1350
rect 131 -1350 165 1350
rect -69 -1446 69 -1412
<< xpolycontact >>
rect -35 884 35 1316
rect -35 -1316 35 -884
<< xpolyres >>
rect -35 -884 35 884
<< locali >>
rect -165 1412 -69 1446
rect 69 1412 165 1446
rect -165 1350 -131 1412
rect 131 1350 165 1412
rect -165 -1412 -131 -1350
rect 131 -1412 165 -1350
rect -165 -1446 -69 -1412
rect 69 -1446 165 -1412
<< viali >>
rect -19 901 19 1298
rect -19 -1298 19 -901
<< metal1 >>
rect -25 1298 25 1310
rect -25 901 -19 1298
rect 19 901 25 1298
rect -25 889 25 901
rect -25 -901 25 -889
rect -25 -1298 -19 -901
rect 19 -1298 25 -901
rect -25 -1310 25 -1298
<< properties >>
string FIXED_BBOX -148 -1429 148 1429
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 9.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 52.504k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
