magic
tech sky130A
magscale 1 2
timestamp 1717527227
<< metal3 >>
rect -986 812 986 840
rect -986 -812 902 812
rect 966 -812 986 812
rect -986 -840 986 -812
<< via3 >>
rect 902 -812 966 812
<< mimcap >>
rect -946 760 654 800
rect -946 -760 -906 760
rect 614 -760 654 760
rect -946 -800 654 -760
<< mimcapcontact >>
rect -906 -760 614 760
<< metal4 >>
rect 886 812 982 828
rect -907 760 615 761
rect -907 -760 -906 760
rect 614 -760 615 760
rect -907 -761 615 -760
rect 886 -812 902 812
rect 966 -812 982 812
rect 886 -828 982 -812
<< properties >>
string FIXED_BBOX -986 -840 694 840
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 8.00 l 8.00 val 134.08 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
