magic
tech sky130A
magscale 1 2
timestamp 1731723950
<< isosubstrate >>
rect 3992 -292617 17571 -279609
<< nwell >>
rect 3668 -279490 17889 -279310
rect 3668 -292646 3908 -279490
rect 17460 -279508 17889 -279490
rect 17709 -285270 17889 -279508
rect 32362 -283550 38526 -283370
rect 32362 -285270 32542 -283550
rect 17709 -285450 32542 -285270
rect 38286 -286171 38526 -283550
rect 38152 -287265 38526 -286171
rect 38286 -292646 38526 -287265
rect 3668 -292890 38526 -292646
<< mvpsubdiff >>
rect 3489 -279177 3549 -279143
rect 17991 -279177 18056 -279143
rect 3489 -279203 3523 -279177
rect 18022 -279198 18056 -279177
rect 18022 -285103 18056 -285071
rect 32195 -283237 32255 -283203
rect 38627 -283237 38687 -283203
rect 32195 -283263 32229 -283237
rect 38653 -283263 38687 -283237
rect 32195 -285103 32229 -285078
rect 18022 -285137 18081 -285103
rect 32163 -285137 32229 -285103
rect 3489 -293013 3523 -292987
rect 38653 -293013 38687 -292987
rect 3489 -293047 3549 -293013
rect 38627 -293047 38687 -293013
<< mvnsubdiff >>
rect 3734 -279410 3794 -279376
rect 17759 -279410 17823 -279376
rect 3734 -279436 3768 -279410
rect 17789 -279441 17823 -279410
rect 32428 -283470 32488 -283436
rect 38400 -283470 38460 -283436
rect 32428 -283496 32462 -283470
rect 17789 -285336 17823 -285296
rect 32428 -285336 32462 -285302
rect 17789 -285370 17857 -285336
rect 32388 -285370 32462 -285336
rect 38426 -283496 38460 -283470
rect 3734 -292790 3768 -292764
rect 38426 -292790 38460 -292764
rect 3734 -292824 3794 -292790
rect 38400 -292824 38460 -292790
<< mvpsubdiffcont >>
rect 3549 -279177 17991 -279143
rect 3489 -292987 3523 -279203
rect 18022 -285071 18056 -279198
rect 32255 -283237 38627 -283203
rect 32195 -285078 32229 -283263
rect 18081 -285137 32163 -285103
rect 38653 -292987 38687 -283263
rect 3549 -293047 38627 -293013
<< mvnsubdiffcont >>
rect 3794 -279410 17759 -279376
rect 3734 -292764 3768 -279436
rect 17789 -285296 17823 -279441
rect 32488 -283470 38400 -283436
rect 32428 -285302 32462 -283496
rect 17857 -285370 32388 -285336
rect 38426 -292764 38460 -283496
rect 3794 -292824 38400 -292790
<< locali >>
rect 3489 -279177 3549 -279143
rect 17991 -279177 18056 -279143
rect 3489 -279198 18056 -279177
rect 3489 -279203 18022 -279198
rect 3523 -279214 18022 -279203
rect 3523 -279260 3551 -279214
rect 3523 -279310 17939 -279260
rect 3523 -279347 3633 -279310
rect 3523 -292843 3540 -279347
rect 3583 -292843 3633 -279347
rect 3734 -279410 3794 -279376
rect 17759 -279410 17823 -279376
rect 3734 -279436 17823 -279410
rect 3768 -279441 17823 -279436
rect 3768 -279446 17789 -279441
rect 3768 -279490 3804 -279446
rect 3768 -279530 17709 -279490
rect 3768 -279548 3895 -279530
rect 3768 -292656 3802 -279548
rect 3844 -292656 3895 -279548
rect 6858 -279717 16036 -279714
rect 6797 -279760 16036 -279717
rect 6797 -279801 7003 -279760
rect 6797 -289021 6865 -279801
rect 6917 -279816 7003 -279801
rect 15989 -279816 16036 -279760
rect 6917 -279903 16036 -279816
rect 6917 -288909 6986 -279903
rect 11271 -280590 12544 -279903
rect 11271 -288849 11530 -280590
rect 12322 -288849 12544 -280590
rect 11271 -288909 12544 -288849
rect 15161 -279908 16036 -279903
rect 15161 -280092 15958 -279908
rect 15161 -280550 15423 -280092
rect 15161 -288909 15216 -280550
rect 6917 -288915 15216 -288909
rect 15268 -281058 15423 -280550
rect 15892 -280998 15958 -280092
rect 16018 -280998 16036 -279908
rect 15892 -281058 16036 -280998
rect 15268 -281202 16036 -281058
rect 15268 -288909 15350 -281202
rect 17669 -285450 17709 -279530
rect 17753 -285296 17789 -279446
rect 17889 -285220 17939 -279310
rect 17985 -285071 18022 -279214
rect 17985 -285103 18056 -285071
rect 32195 -283237 32255 -283203
rect 38627 -283237 38687 -283203
rect 32195 -283263 38687 -283237
rect 32229 -283274 38653 -283263
rect 32229 -283320 32257 -283274
rect 38510 -283306 38653 -283274
rect 38510 -283320 38595 -283306
rect 32229 -283370 38595 -283320
rect 32229 -283407 32362 -283370
rect 32229 -285078 32266 -283407
rect 32195 -285103 32266 -285078
rect 17985 -285137 18081 -285103
rect 32163 -285137 32266 -285103
rect 17985 -285174 32266 -285137
rect 32312 -285220 32362 -283407
rect 17889 -285270 32362 -285220
rect 32428 -283470 32488 -283436
rect 38400 -283470 38460 -283436
rect 32428 -283496 38460 -283470
rect 17753 -285336 17823 -285296
rect 32462 -283506 38426 -283496
rect 32462 -283550 32498 -283506
rect 38319 -283525 38426 -283506
rect 38319 -283550 38363 -283525
rect 32462 -283590 38363 -283550
rect 32462 -283608 32582 -283590
rect 32462 -285302 32498 -283608
rect 32428 -285336 32498 -285302
rect 17753 -285370 17857 -285336
rect 32388 -285370 32498 -285336
rect 17753 -285406 32498 -285370
rect 32542 -285450 32582 -283608
rect 17669 -285490 32582 -285450
rect 15268 -288915 15690 -288909
rect 6917 -288987 15690 -288915
rect 6917 -289021 6984 -288987
rect 6797 -289047 6984 -289021
rect 9475 -289013 15690 -288987
rect 9475 -289047 13305 -289013
rect 6797 -289062 13305 -289047
rect 15607 -289062 15690 -289013
rect 6797 -289098 15690 -289062
rect 9850 -289841 10066 -289098
rect 10476 -289099 13244 -289098
rect 10645 -289165 13244 -289099
rect 10645 -289218 10720 -289165
rect 13220 -289218 13244 -289165
rect 10645 -289355 13244 -289218
rect 10645 -289362 11046 -289355
rect 10645 -289841 10757 -289362
rect 9850 -290003 10757 -289841
rect 9850 -290591 9997 -290003
rect 10476 -290591 10757 -290003
rect 9850 -290755 10757 -290591
rect 9850 -290757 9997 -290755
rect 3768 -292692 3895 -292656
rect 38324 -292692 38363 -283590
rect 3768 -292732 38363 -292692
rect 3768 -292764 3821 -292732
rect 3734 -292769 3821 -292764
rect 38284 -292746 38363 -292732
rect 38402 -292746 38426 -283525
rect 38284 -292764 38426 -292746
rect 38284 -292769 38460 -292764
rect 3734 -292790 38460 -292769
rect 3734 -292824 3794 -292790
rect 38400 -292824 38460 -292790
rect 3523 -292877 3633 -292843
rect 38553 -292873 38595 -283370
rect 38634 -292873 38653 -283306
rect 38553 -292877 38653 -292873
rect 3523 -292942 38653 -292877
rect 3523 -292981 3593 -292942
rect 38616 -292981 38653 -292942
rect 3523 -292987 38653 -292981
rect 3489 -293013 38687 -292987
rect 3489 -293047 3549 -293013
rect 38627 -293047 38687 -293013
<< viali >>
rect 3551 -279260 17985 -279214
rect 3540 -292843 3583 -279347
rect 3804 -279490 17753 -279446
rect 3802 -292656 3844 -279548
rect 6865 -289021 6917 -279801
rect 7003 -279816 15989 -279760
rect 15216 -288915 15268 -280550
rect 15958 -280998 16018 -279908
rect 17709 -285406 17753 -279490
rect 17939 -285174 17985 -279260
rect 32257 -283320 38510 -283274
rect 32266 -285174 32312 -283407
rect 17939 -285220 32312 -285174
rect 32498 -283550 38319 -283506
rect 32498 -285406 32542 -283608
rect 17709 -285450 32542 -285406
rect 6984 -289047 9475 -288987
rect 13305 -289062 15607 -289013
rect 10720 -289218 13220 -289165
rect 3821 -292769 38284 -292732
rect 38363 -292746 38402 -283525
rect 38595 -292873 38634 -283306
rect 3593 -292981 38616 -292942
<< metal1 >>
rect 3493 -279214 18049 -279150
rect 3493 -279260 3551 -279214
rect 3493 -279302 17939 -279260
rect 3502 -279347 3612 -279302
rect 3502 -292843 3540 -279347
rect 3583 -292843 3612 -279347
rect 3756 -279436 17806 -279393
rect 3756 -279446 6368 -279436
rect 3756 -279490 3804 -279446
rect 3756 -279508 6368 -279490
rect 17754 -279508 17806 -279436
rect 3756 -279519 17709 -279508
rect 3756 -279548 3877 -279519
rect 3756 -289178 3802 -279548
rect 3844 -289178 3877 -279548
rect 6800 -279715 7018 -279713
rect 6800 -279760 16046 -279715
rect 6800 -279801 7003 -279760
rect 6800 -279840 6865 -279801
rect 6917 -279816 7003 -279801
rect 15989 -279816 16046 -279760
rect 6800 -288899 6832 -279840
rect 6917 -279894 16046 -279816
rect 6917 -279997 7018 -279894
rect 15145 -279897 16046 -279894
rect 15947 -279908 16046 -279897
rect 6917 -280429 7181 -279997
rect 7277 -280429 7513 -279997
rect 7609 -280429 7845 -279997
rect 7941 -280429 8177 -279997
rect 8273 -280429 8509 -279997
rect 8605 -280429 8841 -279997
rect 8937 -280429 9173 -279997
rect 9269 -280429 9505 -279997
rect 9601 -280429 9837 -279997
rect 9933 -280429 10169 -279997
rect 10265 -280429 10501 -279997
rect 10597 -280429 10833 -279997
rect 10929 -280429 11165 -279997
rect 12634 -280429 12872 -279996
rect 12968 -280429 13206 -279996
rect 13302 -280429 13540 -279996
rect 13636 -280429 13874 -279996
rect 13970 -280429 14208 -279996
rect 14304 -280429 14542 -279996
rect 14638 -280429 14876 -279996
rect 6800 -289021 6865 -288899
rect 6917 -288907 7018 -280429
rect 14983 -280431 15545 -279996
rect 15579 -280228 15758 -280184
rect 15648 -280500 15692 -280228
rect 15145 -280550 15350 -280501
rect 15579 -280542 15746 -280500
rect 11633 -281148 11869 -280715
rect 11964 -281149 12200 -280716
rect 11798 -288225 12340 -288052
rect 7111 -288829 7347 -288397
rect 7443 -288829 7679 -288397
rect 7775 -288829 8011 -288397
rect 8107 -288829 8343 -288397
rect 8439 -288829 8675 -288397
rect 8771 -288829 9007 -288397
rect 9103 -288829 9339 -288397
rect 9435 -288829 9671 -288397
rect 9767 -288829 10003 -288397
rect 10099 -288829 10335 -288397
rect 10431 -288829 10667 -288397
rect 10763 -288829 10999 -288397
rect 11093 -288747 11702 -288397
rect 11388 -288868 11435 -288747
rect 11798 -288748 11869 -288225
rect 6917 -288976 9555 -288907
rect 6917 -289021 6972 -288976
rect 6800 -289052 6972 -289021
rect 9520 -289052 9555 -288976
rect 6800 -289094 9555 -289052
rect 10088 -288915 11435 -288868
rect 7406 -289096 8379 -289094
rect 3756 -289467 3772 -289178
rect 3870 -289467 3877 -289178
rect 10088 -289262 10135 -288915
rect 11965 -288963 12035 -288316
rect 12130 -288394 12340 -288225
rect 12130 -288451 12707 -288394
rect 12135 -288659 12707 -288451
rect 12131 -288748 12707 -288659
rect 10289 -289011 12035 -288963
rect 3756 -292656 3802 -289467
rect 3844 -292656 3877 -289467
rect 10289 -289596 10337 -289011
rect 12382 -289053 12430 -288748
rect 12800 -288829 13038 -288396
rect 13134 -288829 13372 -288396
rect 13468 -288829 13706 -288396
rect 13802 -288829 14040 -288396
rect 14136 -288829 14374 -288396
rect 14470 -288829 14708 -288396
rect 14804 -288829 15042 -288396
rect 15145 -288915 15216 -280550
rect 15268 -288915 15350 -280550
rect 15648 -280608 15692 -280542
rect 15579 -280650 15746 -280608
rect 15417 -281128 15532 -280696
rect 15648 -280922 15692 -280650
rect 15791 -280880 15885 -280270
rect 15579 -280989 15746 -280922
rect 15648 -281128 15692 -280989
rect 15947 -280998 15958 -279908
rect 16018 -280998 16046 -279908
rect 15947 -281023 16046 -280998
rect 15417 -281376 16312 -281128
rect 16605 -281376 16619 -281128
rect 17680 -285450 17709 -279519
rect 17753 -285353 17806 -279508
rect 17897 -285220 17939 -279302
rect 17985 -285110 18049 -279214
rect 32199 -283274 38674 -283210
rect 32199 -283320 32257 -283274
rect 38510 -283306 38674 -283274
rect 38510 -283320 38595 -283306
rect 32199 -283362 38595 -283320
rect 32202 -283407 32354 -283362
rect 32202 -285110 32266 -283407
rect 17985 -285174 32266 -285110
rect 32312 -285220 32354 -283407
rect 17897 -285262 32354 -285220
rect 32445 -283457 38440 -283453
rect 32445 -283506 38447 -283457
rect 32445 -283550 32498 -283506
rect 38319 -283525 38447 -283506
rect 38319 -283550 38363 -283525
rect 32445 -283579 38363 -283550
rect 32445 -283608 32571 -283579
rect 32445 -285353 32498 -283608
rect 17753 -285406 32498 -285353
rect 32542 -285450 32571 -283608
rect 17680 -285479 32571 -285450
rect 15145 -288972 15350 -288915
rect 10484 -289101 12430 -289053
rect 12582 -288976 15663 -288972
rect 12582 -289013 13403 -288976
rect 15496 -289013 15663 -288976
rect 12582 -289062 13305 -289013
rect 15607 -289062 15663 -289013
rect 12582 -289092 15663 -289062
rect 10484 -289210 10532 -289101
rect 12582 -289140 13263 -289092
rect 10686 -289165 13263 -289140
rect 10686 -289218 10720 -289165
rect 13220 -289192 13263 -289165
rect 13220 -289218 13240 -289192
rect 10686 -289348 13240 -289218
rect 11027 -289355 13240 -289348
rect 10048 -290201 10114 -290096
rect 10048 -290408 10132 -290201
rect 10204 -290876 10246 -290137
rect 10353 -290400 10417 -290083
rect 17538 -290701 17586 -289045
rect 16990 -290749 17586 -290701
rect 3756 -292703 3877 -292656
rect 16806 -292530 16892 -292263
rect 16806 -292555 16982 -292530
rect 16806 -292610 17821 -292555
rect 16806 -292611 23772 -292610
rect 16806 -292673 17821 -292611
rect 38334 -292703 38363 -283579
rect 3756 -292732 38363 -292703
rect 3756 -292769 3821 -292732
rect 38284 -292746 38363 -292732
rect 38402 -292746 38447 -283525
rect 38284 -292769 38447 -292746
rect 3756 -292802 38447 -292769
rect 3756 -292805 38380 -292802
rect 3758 -292809 38380 -292805
rect 3502 -292902 3612 -292843
rect 38562 -292873 38595 -283362
rect 38634 -283362 38674 -283306
rect 38634 -292873 38672 -283362
rect 38562 -292902 38672 -292873
rect 3502 -292927 38672 -292902
rect 3502 -292942 17403 -292927
rect 24818 -292942 38672 -292927
rect 3502 -292981 3593 -292942
rect 38616 -292981 38672 -292942
rect 3502 -293001 17403 -292981
rect 24818 -293001 38672 -292981
rect 3502 -293032 38672 -293001
rect 38562 -293043 38672 -293032
<< via1 >>
rect 6368 -279446 17754 -279436
rect 6368 -279490 17753 -279446
rect 6368 -279508 17709 -279490
rect 17709 -279508 17753 -279490
rect 17753 -279508 17754 -279446
rect 6832 -288899 6865 -279840
rect 6865 -288899 6908 -279840
rect 6972 -288987 9520 -288976
rect 6972 -289047 6984 -288987
rect 6984 -289047 9475 -288987
rect 9475 -289047 9520 -288987
rect 6972 -289052 9520 -289047
rect 3772 -289467 3802 -289178
rect 3802 -289467 3844 -289178
rect 3844 -289467 3870 -289178
rect 16312 -281376 16605 -281128
rect 13403 -289013 15496 -288976
rect 13403 -289041 15496 -289013
rect 16786 -289428 17380 -289293
rect 5791 -292476 9241 -292342
rect 12676 -292483 16558 -292395
rect 17403 -292942 24818 -292927
rect 17403 -292981 24818 -292942
rect 17403 -293001 24818 -292981
<< metal2 >>
rect 6314 -279436 17834 -279397
rect 6314 -279497 6368 -279436
rect 6312 -279508 6368 -279497
rect 17754 -279508 17834 -279436
rect 6312 -279652 17834 -279508
rect 6312 -279660 6605 -279652
rect 6705 -279840 6971 -279763
rect 6705 -288899 6832 -279840
rect 6908 -288806 6971 -279840
rect 16312 -281128 16605 -279652
rect 16312 -284876 16605 -281376
rect 39229 -284155 39429 -284118
rect 37892 -284274 39429 -284155
rect 39229 -284318 39429 -284274
rect 24237 -284876 24891 -284875
rect 16312 -285327 24891 -284876
rect 39229 -284905 39429 -284868
rect 37892 -285024 39429 -284905
rect 39229 -285068 39429 -285024
rect 6908 -288899 15690 -288806
rect 6705 -288976 15690 -288899
rect 6705 -289052 6972 -288976
rect 9520 -289041 13403 -288976
rect 15496 -289041 15690 -288976
rect 9520 -289052 15690 -289041
rect 6705 -289072 15690 -289052
rect 3464 -289178 4428 -289169
rect 3464 -289467 3772 -289178
rect 3870 -289467 4428 -289178
rect 16312 -289183 16605 -285327
rect 24237 -285850 24891 -285327
rect 24238 -286408 24891 -285850
rect 3464 -289479 4428 -289467
rect 15582 -289476 16605 -289183
rect 16747 -288187 17828 -287923
rect 16747 -289293 17438 -288187
rect 17564 -289223 17676 -289023
rect 39296 -289256 39496 -289188
rect 16747 -289428 16786 -289293
rect 17380 -289428 17438 -289293
rect 38044 -289340 39496 -289256
rect 39296 -289388 39496 -289340
rect 16747 -289466 17438 -289428
rect 10326 -290222 10378 -289565
rect 37864 -290005 39496 -289913
rect 35038 -290006 39496 -290005
rect 35038 -290381 39497 -290006
rect 37864 -290493 39496 -290381
rect 39301 -290786 39501 -290729
rect 37952 -290871 39501 -290786
rect 37952 -291076 38037 -290871
rect 39301 -290929 39501 -290871
rect 4462 -292342 9298 -292313
rect 4462 -292476 5791 -292342
rect 9241 -292476 9298 -292342
rect 4462 -292805 9298 -292476
rect 12630 -292395 16597 -292360
rect 12630 -292483 12676 -292395
rect 16558 -292483 16597 -292395
rect 12630 -292805 16597 -292483
rect 4462 -292806 16600 -292805
rect 3564 -293345 16600 -292806
rect 4462 -293347 16600 -293345
rect 17324 -292927 17872 -292805
rect 17324 -293001 17403 -292927
rect 17324 -293003 17872 -293001
rect 17324 -293338 24877 -293003
rect 17324 -293347 17872 -293338
<< metal3 >>
rect 32079 -284981 32641 -284194
<< metal4 >>
rect 32079 -284981 32641 -284194
<< metal5 >>
rect 32079 -284981 32641 -284194
use por_via_2cut  por_via_2cut_0
timestamp 1718283729
transform 0 1 18285 -1 0 -274010
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_2
timestamp 1718283729
transform -1 0 26472 0 -1 -297476
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_4
timestamp 1718283729
transform 0 1 17981 -1 0 -274025
box 16088 -7932 16222 -7868
use por_via_4cut  por_via_4cut_18
timestamp 1718283729
transform 0 -1 9666 1 0 -305206
box 15948 -7932 16222 -7868
use sky130_fd_pr__res_xhigh_po_0p35_WGPHGK  R1 paramcells
timestamp 1731359787
transform 1 0 9138 0 1 -284414
box -2193 -4582 2193 4582
use sky130_fd_pr__res_xhigh_po_0p35_PXB2PH  R10 paramcells
timestamp 1731450921
transform 1 0 11917 0 1 -284732
box -450 -4182 450 4182
use sky130_fd_pr__res_xhigh_po_0p35_MNWQZD  R12 paramcells
timestamp 1731359787
transform 1 0 13835 0 1 -284412
box -1363 -4582 1363 4582
use sky130_fd_pr__nfet_05v0_nvt_FPTPS4  sky130_fd_pr__nfet_05v0_nvt_FPTPS4_0 paramcells
timestamp 1731450921
transform 1 0 10231 0 1 -290301
box -318 -358 318 358
use comparator_final  x1
timestamp 1731723950
transform 1 0 6296 0 1 -286728
box -1988 -5804 11208 -2441
use delayPulse_final  x2
timestamp 1731723950
transform 1 0 1055 0 1 -2959
box 1311 -297437 38614 -274935
use sky130_fd_pr__nfet_05v0_nvt_CZFQWY  XM2 paramcells
timestamp 1726591550
transform 1 0 15668 0 1 -280576
box -318 -567 318 567
<< labels >>
flabel metal2 39296 -289388 39496 -289188 0 FreeSans 256 0 0 0 porb
port 5 nsew
flabel metal2 39301 -290929 39501 -290729 0 FreeSans 256 0 0 0 por
port 1 nsew
flabel metal2 24555 -293294 24755 -293094 0 FreeSans 256 0 0 0 dvss
port 6 nsew
flabel metal2 39292 -290256 39492 -290056 0 FreeSans 256 0 0 0 dvdd
port 4 nsew
flabel metal2 3491 -289455 3691 -289255 0 FreeSans 256 0 0 0 avdd
port 3 nsew
flabel metal2 3612 -293264 3812 -293064 0 FreeSans 256 0 0 0 avss
port 2 nsew
flabel metal2 39229 -285068 39429 -284868 0 FreeSans 256 0 0 0 porb_h[1]
port 8 nsew
flabel metal2 39229 -284318 39429 -284118 0 FreeSans 256 0 0 0 porb_h[0]
port 7 nsew
<< end >>
