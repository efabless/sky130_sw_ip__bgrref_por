magic
tech sky130A
magscale 1 2
timestamp 1718283729
<< metal3 >>
rect -4192 18154 -566 18182
rect -4192 14930 -650 18154
rect -586 14930 -566 18154
rect -4192 14902 -566 14930
rect 120 18154 3746 18182
rect 120 14930 3662 18154
rect 3726 14930 3746 18154
rect 120 14902 3746 14930
rect -4192 14556 -566 14584
rect -4192 11332 -650 14556
rect -586 11332 -566 14556
rect -4192 11304 -566 11332
rect 120 14556 3746 14584
rect 120 11332 3662 14556
rect 3726 11332 3746 14556
rect 120 11304 3746 11332
rect -4192 10958 -566 10986
rect -4192 7734 -650 10958
rect -586 7734 -566 10958
rect -4192 7706 -566 7734
rect 120 10958 3746 10986
rect 120 7734 3662 10958
rect 3726 7734 3746 10958
rect 120 7706 3746 7734
rect -4192 7360 -566 7388
rect -4192 4136 -650 7360
rect -586 4136 -566 7360
rect -4192 4108 -566 4136
rect 120 7360 3746 7388
rect 120 4136 3662 7360
rect 3726 4136 3746 7360
rect 120 4108 3746 4136
rect -4192 3762 -566 3790
rect -4192 538 -650 3762
rect -586 538 -566 3762
rect -4192 510 -566 538
rect 120 3762 3746 3790
rect 120 538 3662 3762
rect 3726 538 3746 3762
rect 120 510 3746 538
rect -4192 164 -566 192
rect -4192 -3060 -650 164
rect -586 -3060 -566 164
rect -4192 -3088 -566 -3060
rect 120 164 3746 192
rect 120 -3060 3662 164
rect 3726 -3060 3746 164
rect 120 -3088 3746 -3060
rect -4192 -3434 -566 -3406
rect -4192 -6658 -650 -3434
rect -586 -6658 -566 -3434
rect -4192 -6686 -566 -6658
rect 120 -3434 3746 -3406
rect 120 -6658 3662 -3434
rect 3726 -6658 3746 -3434
rect 120 -6686 3746 -6658
rect -4192 -7032 -566 -7004
rect -4192 -10256 -650 -7032
rect -586 -10256 -566 -7032
rect -4192 -10284 -566 -10256
rect 120 -7032 3746 -7004
rect 120 -10256 3662 -7032
rect 3726 -10256 3746 -7032
rect 120 -10284 3746 -10256
rect -4192 -10630 -566 -10602
rect -4192 -13854 -650 -10630
rect -586 -13854 -566 -10630
rect -4192 -13882 -566 -13854
rect 120 -10630 3746 -10602
rect 120 -13854 3662 -10630
rect 3726 -13854 3746 -10630
rect 120 -13882 3746 -13854
rect -4192 -14228 -566 -14200
rect -4192 -17452 -650 -14228
rect -586 -17452 -566 -14228
rect -4192 -17480 -566 -17452
rect 120 -14228 3746 -14200
rect 120 -17452 3662 -14228
rect 3726 -17452 3746 -14228
rect 120 -17480 3746 -17452
<< via3 >>
rect -650 14930 -586 18154
rect 3662 14930 3726 18154
rect -650 11332 -586 14556
rect 3662 11332 3726 14556
rect -650 7734 -586 10958
rect 3662 7734 3726 10958
rect -650 4136 -586 7360
rect 3662 4136 3726 7360
rect -650 538 -586 3762
rect 3662 538 3726 3762
rect -650 -3060 -586 164
rect 3662 -3060 3726 164
rect -650 -6658 -586 -3434
rect 3662 -6658 3726 -3434
rect -650 -10256 -586 -7032
rect 3662 -10256 3726 -7032
rect -650 -13854 -586 -10630
rect 3662 -13854 3726 -10630
rect -650 -17452 -586 -14228
rect 3662 -17452 3726 -14228
<< mimcap >>
rect -4152 18102 -952 18142
rect -4152 14982 -4112 18102
rect -992 14982 -952 18102
rect -4152 14942 -952 14982
rect 160 18102 3360 18142
rect 160 14982 200 18102
rect 3320 14982 3360 18102
rect 160 14942 3360 14982
rect -4152 14504 -952 14544
rect -4152 11384 -4112 14504
rect -992 11384 -952 14504
rect -4152 11344 -952 11384
rect 160 14504 3360 14544
rect 160 11384 200 14504
rect 3320 11384 3360 14504
rect 160 11344 3360 11384
rect -4152 10906 -952 10946
rect -4152 7786 -4112 10906
rect -992 7786 -952 10906
rect -4152 7746 -952 7786
rect 160 10906 3360 10946
rect 160 7786 200 10906
rect 3320 7786 3360 10906
rect 160 7746 3360 7786
rect -4152 7308 -952 7348
rect -4152 4188 -4112 7308
rect -992 4188 -952 7308
rect -4152 4148 -952 4188
rect 160 7308 3360 7348
rect 160 4188 200 7308
rect 3320 4188 3360 7308
rect 160 4148 3360 4188
rect -4152 3710 -952 3750
rect -4152 590 -4112 3710
rect -992 590 -952 3710
rect -4152 550 -952 590
rect 160 3710 3360 3750
rect 160 590 200 3710
rect 3320 590 3360 3710
rect 160 550 3360 590
rect -4152 112 -952 152
rect -4152 -3008 -4112 112
rect -992 -3008 -952 112
rect -4152 -3048 -952 -3008
rect 160 112 3360 152
rect 160 -3008 200 112
rect 3320 -3008 3360 112
rect 160 -3048 3360 -3008
rect -4152 -3486 -952 -3446
rect -4152 -6606 -4112 -3486
rect -992 -6606 -952 -3486
rect -4152 -6646 -952 -6606
rect 160 -3486 3360 -3446
rect 160 -6606 200 -3486
rect 3320 -6606 3360 -3486
rect 160 -6646 3360 -6606
rect -4152 -7084 -952 -7044
rect -4152 -10204 -4112 -7084
rect -992 -10204 -952 -7084
rect -4152 -10244 -952 -10204
rect 160 -7084 3360 -7044
rect 160 -10204 200 -7084
rect 3320 -10204 3360 -7084
rect 160 -10244 3360 -10204
rect -4152 -10682 -952 -10642
rect -4152 -13802 -4112 -10682
rect -992 -13802 -952 -10682
rect -4152 -13842 -952 -13802
rect 160 -10682 3360 -10642
rect 160 -13802 200 -10682
rect 3320 -13802 3360 -10682
rect 160 -13842 3360 -13802
rect -4152 -14280 -952 -14240
rect -4152 -17400 -4112 -14280
rect -992 -17400 -952 -14280
rect -4152 -17440 -952 -17400
rect 160 -14280 3360 -14240
rect 160 -17400 200 -14280
rect 3320 -17400 3360 -14280
rect 160 -17440 3360 -17400
<< mimcapcontact >>
rect -4112 14982 -992 18102
rect 200 14982 3320 18102
rect -4112 11384 -992 14504
rect 200 11384 3320 14504
rect -4112 7786 -992 10906
rect 200 7786 3320 10906
rect -4112 4188 -992 7308
rect 200 4188 3320 7308
rect -4112 590 -992 3710
rect 200 590 3320 3710
rect -4112 -3008 -992 112
rect 200 -3008 3320 112
rect -4112 -6606 -992 -3486
rect 200 -6606 3320 -3486
rect -4112 -10204 -992 -7084
rect 200 -10204 3320 -7084
rect -4112 -13802 -992 -10682
rect 200 -13802 3320 -10682
rect -4112 -17400 -992 -14280
rect 200 -17400 3320 -14280
<< metal4 >>
rect -2604 18103 -2500 18302
rect -670 18154 -566 18302
rect -4113 18102 -991 18103
rect -4113 14982 -4112 18102
rect -992 14982 -991 18102
rect -4113 14981 -991 14982
rect -2604 14505 -2500 14981
rect -670 14930 -650 18154
rect -586 14930 -566 18154
rect 1708 18103 1812 18302
rect 3642 18154 3746 18302
rect 199 18102 3321 18103
rect 199 14982 200 18102
rect 3320 14982 3321 18102
rect 199 14981 3321 14982
rect -670 14556 -566 14930
rect -4113 14504 -991 14505
rect -4113 11384 -4112 14504
rect -992 11384 -991 14504
rect -4113 11383 -991 11384
rect -2604 10907 -2500 11383
rect -670 11332 -650 14556
rect -586 11332 -566 14556
rect 1708 14505 1812 14981
rect 3642 14930 3662 18154
rect 3726 14930 3746 18154
rect 3642 14556 3746 14930
rect 199 14504 3321 14505
rect 199 11384 200 14504
rect 3320 11384 3321 14504
rect 199 11383 3321 11384
rect -670 10958 -566 11332
rect -4113 10906 -991 10907
rect -4113 7786 -4112 10906
rect -992 7786 -991 10906
rect -4113 7785 -991 7786
rect -2604 7309 -2500 7785
rect -670 7734 -650 10958
rect -586 7734 -566 10958
rect 1708 10907 1812 11383
rect 3642 11332 3662 14556
rect 3726 11332 3746 14556
rect 3642 10958 3746 11332
rect 199 10906 3321 10907
rect 199 7786 200 10906
rect 3320 7786 3321 10906
rect 199 7785 3321 7786
rect -670 7360 -566 7734
rect -4113 7308 -991 7309
rect -4113 4188 -4112 7308
rect -992 4188 -991 7308
rect -4113 4187 -991 4188
rect -2604 3711 -2500 4187
rect -670 4136 -650 7360
rect -586 4136 -566 7360
rect 1708 7309 1812 7785
rect 3642 7734 3662 10958
rect 3726 7734 3746 10958
rect 3642 7360 3746 7734
rect 199 7308 3321 7309
rect 199 4188 200 7308
rect 3320 4188 3321 7308
rect 199 4187 3321 4188
rect -670 3762 -566 4136
rect -4113 3710 -991 3711
rect -4113 590 -4112 3710
rect -992 590 -991 3710
rect -4113 589 -991 590
rect -2604 113 -2500 589
rect -670 538 -650 3762
rect -586 538 -566 3762
rect 1708 3711 1812 4187
rect 3642 4136 3662 7360
rect 3726 4136 3746 7360
rect 3642 3762 3746 4136
rect 199 3710 3321 3711
rect 199 590 200 3710
rect 3320 590 3321 3710
rect 199 589 3321 590
rect -670 164 -566 538
rect -4113 112 -991 113
rect -4113 -3008 -4112 112
rect -992 -3008 -991 112
rect -4113 -3009 -991 -3008
rect -2604 -3485 -2500 -3009
rect -670 -3060 -650 164
rect -586 -3060 -566 164
rect 1708 113 1812 589
rect 3642 538 3662 3762
rect 3726 538 3746 3762
rect 3642 164 3746 538
rect 199 112 3321 113
rect 199 -3008 200 112
rect 3320 -3008 3321 112
rect 199 -3009 3321 -3008
rect -670 -3434 -566 -3060
rect -4113 -3486 -991 -3485
rect -4113 -6606 -4112 -3486
rect -992 -6606 -991 -3486
rect -4113 -6607 -991 -6606
rect -2604 -7083 -2500 -6607
rect -670 -6658 -650 -3434
rect -586 -6658 -566 -3434
rect 1708 -3485 1812 -3009
rect 3642 -3060 3662 164
rect 3726 -3060 3746 164
rect 3642 -3434 3746 -3060
rect 199 -3486 3321 -3485
rect 199 -6606 200 -3486
rect 3320 -6606 3321 -3486
rect 199 -6607 3321 -6606
rect -670 -7032 -566 -6658
rect -4113 -7084 -991 -7083
rect -4113 -10204 -4112 -7084
rect -992 -10204 -991 -7084
rect -4113 -10205 -991 -10204
rect -2604 -10681 -2500 -10205
rect -670 -10256 -650 -7032
rect -586 -10256 -566 -7032
rect 1708 -7083 1812 -6607
rect 3642 -6658 3662 -3434
rect 3726 -6658 3746 -3434
rect 3642 -7032 3746 -6658
rect 199 -7084 3321 -7083
rect 199 -10204 200 -7084
rect 3320 -10204 3321 -7084
rect 199 -10205 3321 -10204
rect -670 -10630 -566 -10256
rect -4113 -10682 -991 -10681
rect -4113 -13802 -4112 -10682
rect -992 -13802 -991 -10682
rect -4113 -13803 -991 -13802
rect -2604 -14279 -2500 -13803
rect -670 -13854 -650 -10630
rect -586 -13854 -566 -10630
rect 1708 -10681 1812 -10205
rect 3642 -10256 3662 -7032
rect 3726 -10256 3746 -7032
rect 3642 -10630 3746 -10256
rect 199 -10682 3321 -10681
rect 199 -13802 200 -10682
rect 3320 -13802 3321 -10682
rect 199 -13803 3321 -13802
rect -670 -14228 -566 -13854
rect -4113 -14280 -991 -14279
rect -4113 -17400 -4112 -14280
rect -992 -17400 -991 -14280
rect -4113 -17401 -991 -17400
rect -2604 -17600 -2500 -17401
rect -670 -17452 -650 -14228
rect -586 -17452 -566 -14228
rect 1708 -14279 1812 -13803
rect 3642 -13854 3662 -10630
rect 3726 -13854 3746 -10630
rect 3642 -14228 3746 -13854
rect 199 -14280 3321 -14279
rect 199 -17400 200 -14280
rect 3320 -17400 3321 -14280
rect 199 -17401 3321 -17400
rect -670 -17600 -566 -17452
rect 1708 -17600 1812 -17401
rect 3642 -17452 3662 -14228
rect 3726 -17452 3746 -14228
rect 3642 -17600 3746 -17452
<< properties >>
string FIXED_BBOX 120 14200 3400 17480
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 16.00 l 16.00 val 524.159 carea 2.00 cperi 0.19 nx 2 ny 10 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
