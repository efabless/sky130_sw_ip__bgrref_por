magic
tech sky130A
magscale 1 2
timestamp 1717363523
<< error_p >>
rect -77 2971 -19 2977
rect -77 2937 -65 2971
rect -77 2931 -19 2937
rect 19 2703 77 2709
rect 19 2669 31 2703
rect 19 2663 77 2669
rect 19 2595 77 2601
rect 19 2561 31 2595
rect 19 2555 77 2561
rect -77 2327 -19 2333
rect -77 2293 -65 2327
rect -77 2287 -19 2293
rect -77 2219 -19 2225
rect -77 2185 -65 2219
rect -77 2179 -19 2185
rect 19 1951 77 1957
rect 19 1917 31 1951
rect 19 1911 77 1917
rect 19 1843 77 1849
rect 19 1809 31 1843
rect 19 1803 77 1809
rect -77 1575 -19 1581
rect -77 1541 -65 1575
rect -77 1535 -19 1541
rect -77 1467 -19 1473
rect -77 1433 -65 1467
rect -77 1427 -19 1433
rect 19 1199 77 1205
rect 19 1165 31 1199
rect 19 1159 77 1165
rect 19 1091 77 1097
rect 19 1057 31 1091
rect 19 1051 77 1057
rect -77 823 -19 829
rect -77 789 -65 823
rect -77 783 -19 789
rect -77 715 -19 721
rect -77 681 -65 715
rect -77 675 -19 681
rect 19 447 77 453
rect 19 413 31 447
rect 19 407 77 413
rect 19 339 77 345
rect 19 305 31 339
rect 19 299 77 305
rect -77 71 -19 77
rect -77 37 -65 71
rect -77 31 -19 37
rect -77 -37 -19 -31
rect -77 -71 -65 -37
rect -77 -77 -19 -71
rect 19 -305 77 -299
rect 19 -339 31 -305
rect 19 -345 77 -339
rect 19 -413 77 -407
rect 19 -447 31 -413
rect 19 -453 77 -447
rect -77 -681 -19 -675
rect -77 -715 -65 -681
rect -77 -721 -19 -715
rect -77 -789 -19 -783
rect -77 -823 -65 -789
rect -77 -829 -19 -823
rect 19 -1057 77 -1051
rect 19 -1091 31 -1057
rect 19 -1097 77 -1091
rect 19 -1165 77 -1159
rect 19 -1199 31 -1165
rect 19 -1205 77 -1199
rect -77 -1433 -19 -1427
rect -77 -1467 -65 -1433
rect -77 -1473 -19 -1467
rect -77 -1541 -19 -1535
rect -77 -1575 -65 -1541
rect -77 -1581 -19 -1575
rect 19 -1809 77 -1803
rect 19 -1843 31 -1809
rect 19 -1849 77 -1843
rect 19 -1917 77 -1911
rect 19 -1951 31 -1917
rect 19 -1957 77 -1951
rect -77 -2185 -19 -2179
rect -77 -2219 -65 -2185
rect -77 -2225 -19 -2219
rect -77 -2293 -19 -2287
rect -77 -2327 -65 -2293
rect -77 -2333 -19 -2327
rect 19 -2561 77 -2555
rect 19 -2595 31 -2561
rect 19 -2601 77 -2595
rect 19 -2669 77 -2663
rect 19 -2703 31 -2669
rect 19 -2709 77 -2703
rect -77 -2937 -19 -2931
rect -77 -2971 -65 -2937
rect -77 -2977 -19 -2971
<< nwell >>
rect -263 -3109 263 3109
<< pmos >>
rect -63 2750 -33 2890
rect 33 2750 63 2890
rect -63 2374 -33 2514
rect 33 2374 63 2514
rect -63 1998 -33 2138
rect 33 1998 63 2138
rect -63 1622 -33 1762
rect 33 1622 63 1762
rect -63 1246 -33 1386
rect 33 1246 63 1386
rect -63 870 -33 1010
rect 33 870 63 1010
rect -63 494 -33 634
rect 33 494 63 634
rect -63 118 -33 258
rect 33 118 63 258
rect -63 -258 -33 -118
rect 33 -258 63 -118
rect -63 -634 -33 -494
rect 33 -634 63 -494
rect -63 -1010 -33 -870
rect 33 -1010 63 -870
rect -63 -1386 -33 -1246
rect 33 -1386 63 -1246
rect -63 -1762 -33 -1622
rect 33 -1762 63 -1622
rect -63 -2138 -33 -1998
rect 33 -2138 63 -1998
rect -63 -2514 -33 -2374
rect 33 -2514 63 -2374
rect -63 -2890 -33 -2750
rect 33 -2890 63 -2750
<< pdiff >>
rect -125 2878 -63 2890
rect -125 2762 -113 2878
rect -79 2762 -63 2878
rect -125 2750 -63 2762
rect -33 2878 33 2890
rect -33 2762 -17 2878
rect 17 2762 33 2878
rect -33 2750 33 2762
rect 63 2878 125 2890
rect 63 2762 79 2878
rect 113 2762 125 2878
rect 63 2750 125 2762
rect -125 2502 -63 2514
rect -125 2386 -113 2502
rect -79 2386 -63 2502
rect -125 2374 -63 2386
rect -33 2502 33 2514
rect -33 2386 -17 2502
rect 17 2386 33 2502
rect -33 2374 33 2386
rect 63 2502 125 2514
rect 63 2386 79 2502
rect 113 2386 125 2502
rect 63 2374 125 2386
rect -125 2126 -63 2138
rect -125 2010 -113 2126
rect -79 2010 -63 2126
rect -125 1998 -63 2010
rect -33 2126 33 2138
rect -33 2010 -17 2126
rect 17 2010 33 2126
rect -33 1998 33 2010
rect 63 2126 125 2138
rect 63 2010 79 2126
rect 113 2010 125 2126
rect 63 1998 125 2010
rect -125 1750 -63 1762
rect -125 1634 -113 1750
rect -79 1634 -63 1750
rect -125 1622 -63 1634
rect -33 1750 33 1762
rect -33 1634 -17 1750
rect 17 1634 33 1750
rect -33 1622 33 1634
rect 63 1750 125 1762
rect 63 1634 79 1750
rect 113 1634 125 1750
rect 63 1622 125 1634
rect -125 1374 -63 1386
rect -125 1258 -113 1374
rect -79 1258 -63 1374
rect -125 1246 -63 1258
rect -33 1374 33 1386
rect -33 1258 -17 1374
rect 17 1258 33 1374
rect -33 1246 33 1258
rect 63 1374 125 1386
rect 63 1258 79 1374
rect 113 1258 125 1374
rect 63 1246 125 1258
rect -125 998 -63 1010
rect -125 882 -113 998
rect -79 882 -63 998
rect -125 870 -63 882
rect -33 998 33 1010
rect -33 882 -17 998
rect 17 882 33 998
rect -33 870 33 882
rect 63 998 125 1010
rect 63 882 79 998
rect 113 882 125 998
rect 63 870 125 882
rect -125 622 -63 634
rect -125 506 -113 622
rect -79 506 -63 622
rect -125 494 -63 506
rect -33 622 33 634
rect -33 506 -17 622
rect 17 506 33 622
rect -33 494 33 506
rect 63 622 125 634
rect 63 506 79 622
rect 113 506 125 622
rect 63 494 125 506
rect -125 246 -63 258
rect -125 130 -113 246
rect -79 130 -63 246
rect -125 118 -63 130
rect -33 246 33 258
rect -33 130 -17 246
rect 17 130 33 246
rect -33 118 33 130
rect 63 246 125 258
rect 63 130 79 246
rect 113 130 125 246
rect 63 118 125 130
rect -125 -130 -63 -118
rect -125 -246 -113 -130
rect -79 -246 -63 -130
rect -125 -258 -63 -246
rect -33 -130 33 -118
rect -33 -246 -17 -130
rect 17 -246 33 -130
rect -33 -258 33 -246
rect 63 -130 125 -118
rect 63 -246 79 -130
rect 113 -246 125 -130
rect 63 -258 125 -246
rect -125 -506 -63 -494
rect -125 -622 -113 -506
rect -79 -622 -63 -506
rect -125 -634 -63 -622
rect -33 -506 33 -494
rect -33 -622 -17 -506
rect 17 -622 33 -506
rect -33 -634 33 -622
rect 63 -506 125 -494
rect 63 -622 79 -506
rect 113 -622 125 -506
rect 63 -634 125 -622
rect -125 -882 -63 -870
rect -125 -998 -113 -882
rect -79 -998 -63 -882
rect -125 -1010 -63 -998
rect -33 -882 33 -870
rect -33 -998 -17 -882
rect 17 -998 33 -882
rect -33 -1010 33 -998
rect 63 -882 125 -870
rect 63 -998 79 -882
rect 113 -998 125 -882
rect 63 -1010 125 -998
rect -125 -1258 -63 -1246
rect -125 -1374 -113 -1258
rect -79 -1374 -63 -1258
rect -125 -1386 -63 -1374
rect -33 -1258 33 -1246
rect -33 -1374 -17 -1258
rect 17 -1374 33 -1258
rect -33 -1386 33 -1374
rect 63 -1258 125 -1246
rect 63 -1374 79 -1258
rect 113 -1374 125 -1258
rect 63 -1386 125 -1374
rect -125 -1634 -63 -1622
rect -125 -1750 -113 -1634
rect -79 -1750 -63 -1634
rect -125 -1762 -63 -1750
rect -33 -1634 33 -1622
rect -33 -1750 -17 -1634
rect 17 -1750 33 -1634
rect -33 -1762 33 -1750
rect 63 -1634 125 -1622
rect 63 -1750 79 -1634
rect 113 -1750 125 -1634
rect 63 -1762 125 -1750
rect -125 -2010 -63 -1998
rect -125 -2126 -113 -2010
rect -79 -2126 -63 -2010
rect -125 -2138 -63 -2126
rect -33 -2010 33 -1998
rect -33 -2126 -17 -2010
rect 17 -2126 33 -2010
rect -33 -2138 33 -2126
rect 63 -2010 125 -1998
rect 63 -2126 79 -2010
rect 113 -2126 125 -2010
rect 63 -2138 125 -2126
rect -125 -2386 -63 -2374
rect -125 -2502 -113 -2386
rect -79 -2502 -63 -2386
rect -125 -2514 -63 -2502
rect -33 -2386 33 -2374
rect -33 -2502 -17 -2386
rect 17 -2502 33 -2386
rect -33 -2514 33 -2502
rect 63 -2386 125 -2374
rect 63 -2502 79 -2386
rect 113 -2502 125 -2386
rect 63 -2514 125 -2502
rect -125 -2762 -63 -2750
rect -125 -2878 -113 -2762
rect -79 -2878 -63 -2762
rect -125 -2890 -63 -2878
rect -33 -2762 33 -2750
rect -33 -2878 -17 -2762
rect 17 -2878 33 -2762
rect -33 -2890 33 -2878
rect 63 -2762 125 -2750
rect 63 -2878 79 -2762
rect 113 -2878 125 -2762
rect 63 -2890 125 -2878
<< pdiffc >>
rect -113 2762 -79 2878
rect -17 2762 17 2878
rect 79 2762 113 2878
rect -113 2386 -79 2502
rect -17 2386 17 2502
rect 79 2386 113 2502
rect -113 2010 -79 2126
rect -17 2010 17 2126
rect 79 2010 113 2126
rect -113 1634 -79 1750
rect -17 1634 17 1750
rect 79 1634 113 1750
rect -113 1258 -79 1374
rect -17 1258 17 1374
rect 79 1258 113 1374
rect -113 882 -79 998
rect -17 882 17 998
rect 79 882 113 998
rect -113 506 -79 622
rect -17 506 17 622
rect 79 506 113 622
rect -113 130 -79 246
rect -17 130 17 246
rect 79 130 113 246
rect -113 -246 -79 -130
rect -17 -246 17 -130
rect 79 -246 113 -130
rect -113 -622 -79 -506
rect -17 -622 17 -506
rect 79 -622 113 -506
rect -113 -998 -79 -882
rect -17 -998 17 -882
rect 79 -998 113 -882
rect -113 -1374 -79 -1258
rect -17 -1374 17 -1258
rect 79 -1374 113 -1258
rect -113 -1750 -79 -1634
rect -17 -1750 17 -1634
rect 79 -1750 113 -1634
rect -113 -2126 -79 -2010
rect -17 -2126 17 -2010
rect 79 -2126 113 -2010
rect -113 -2502 -79 -2386
rect -17 -2502 17 -2386
rect 79 -2502 113 -2386
rect -113 -2878 -79 -2762
rect -17 -2878 17 -2762
rect 79 -2878 113 -2762
<< nsubdiff >>
rect -227 3039 -131 3073
rect 131 3039 227 3073
rect -227 2977 -193 3039
rect 193 2977 227 3039
rect -227 -3039 -193 -2977
rect 193 -3039 227 -2977
rect -227 -3073 -131 -3039
rect 131 -3073 227 -3039
<< nsubdiffcont >>
rect -131 3039 131 3073
rect -227 -2977 -193 2977
rect 193 -2977 227 2977
rect -131 -3073 131 -3039
<< poly >>
rect -81 2971 -15 2987
rect -81 2937 -65 2971
rect -31 2937 -15 2971
rect -81 2921 -15 2937
rect -63 2890 -33 2921
rect 33 2890 63 2916
rect -63 2724 -33 2750
rect 33 2719 63 2750
rect 15 2703 81 2719
rect 15 2669 31 2703
rect 65 2669 81 2703
rect 15 2653 81 2669
rect 15 2595 81 2611
rect 15 2561 31 2595
rect 65 2561 81 2595
rect 15 2545 81 2561
rect -63 2514 -33 2540
rect 33 2514 63 2545
rect -63 2343 -33 2374
rect 33 2348 63 2374
rect -81 2327 -15 2343
rect -81 2293 -65 2327
rect -31 2293 -15 2327
rect -81 2277 -15 2293
rect -81 2219 -15 2235
rect -81 2185 -65 2219
rect -31 2185 -15 2219
rect -81 2169 -15 2185
rect -63 2138 -33 2169
rect 33 2138 63 2164
rect -63 1972 -33 1998
rect 33 1967 63 1998
rect 15 1951 81 1967
rect 15 1917 31 1951
rect 65 1917 81 1951
rect 15 1901 81 1917
rect 15 1843 81 1859
rect 15 1809 31 1843
rect 65 1809 81 1843
rect 15 1793 81 1809
rect -63 1762 -33 1788
rect 33 1762 63 1793
rect -63 1591 -33 1622
rect 33 1596 63 1622
rect -81 1575 -15 1591
rect -81 1541 -65 1575
rect -31 1541 -15 1575
rect -81 1525 -15 1541
rect -81 1467 -15 1483
rect -81 1433 -65 1467
rect -31 1433 -15 1467
rect -81 1417 -15 1433
rect -63 1386 -33 1417
rect 33 1386 63 1412
rect -63 1220 -33 1246
rect 33 1215 63 1246
rect 15 1199 81 1215
rect 15 1165 31 1199
rect 65 1165 81 1199
rect 15 1149 81 1165
rect 15 1091 81 1107
rect 15 1057 31 1091
rect 65 1057 81 1091
rect 15 1041 81 1057
rect -63 1010 -33 1036
rect 33 1010 63 1041
rect -63 839 -33 870
rect 33 844 63 870
rect -81 823 -15 839
rect -81 789 -65 823
rect -31 789 -15 823
rect -81 773 -15 789
rect -81 715 -15 731
rect -81 681 -65 715
rect -31 681 -15 715
rect -81 665 -15 681
rect -63 634 -33 665
rect 33 634 63 660
rect -63 468 -33 494
rect 33 463 63 494
rect 15 447 81 463
rect 15 413 31 447
rect 65 413 81 447
rect 15 397 81 413
rect 15 339 81 355
rect 15 305 31 339
rect 65 305 81 339
rect 15 289 81 305
rect -63 258 -33 284
rect 33 258 63 289
rect -63 87 -33 118
rect 33 92 63 118
rect -81 71 -15 87
rect -81 37 -65 71
rect -31 37 -15 71
rect -81 21 -15 37
rect -81 -37 -15 -21
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect -81 -87 -15 -71
rect -63 -118 -33 -87
rect 33 -118 63 -92
rect -63 -284 -33 -258
rect 33 -289 63 -258
rect 15 -305 81 -289
rect 15 -339 31 -305
rect 65 -339 81 -305
rect 15 -355 81 -339
rect 15 -413 81 -397
rect 15 -447 31 -413
rect 65 -447 81 -413
rect 15 -463 81 -447
rect -63 -494 -33 -468
rect 33 -494 63 -463
rect -63 -665 -33 -634
rect 33 -660 63 -634
rect -81 -681 -15 -665
rect -81 -715 -65 -681
rect -31 -715 -15 -681
rect -81 -731 -15 -715
rect -81 -789 -15 -773
rect -81 -823 -65 -789
rect -31 -823 -15 -789
rect -81 -839 -15 -823
rect -63 -870 -33 -839
rect 33 -870 63 -844
rect -63 -1036 -33 -1010
rect 33 -1041 63 -1010
rect 15 -1057 81 -1041
rect 15 -1091 31 -1057
rect 65 -1091 81 -1057
rect 15 -1107 81 -1091
rect 15 -1165 81 -1149
rect 15 -1199 31 -1165
rect 65 -1199 81 -1165
rect 15 -1215 81 -1199
rect -63 -1246 -33 -1220
rect 33 -1246 63 -1215
rect -63 -1417 -33 -1386
rect 33 -1412 63 -1386
rect -81 -1433 -15 -1417
rect -81 -1467 -65 -1433
rect -31 -1467 -15 -1433
rect -81 -1483 -15 -1467
rect -81 -1541 -15 -1525
rect -81 -1575 -65 -1541
rect -31 -1575 -15 -1541
rect -81 -1591 -15 -1575
rect -63 -1622 -33 -1591
rect 33 -1622 63 -1596
rect -63 -1788 -33 -1762
rect 33 -1793 63 -1762
rect 15 -1809 81 -1793
rect 15 -1843 31 -1809
rect 65 -1843 81 -1809
rect 15 -1859 81 -1843
rect 15 -1917 81 -1901
rect 15 -1951 31 -1917
rect 65 -1951 81 -1917
rect 15 -1967 81 -1951
rect -63 -1998 -33 -1972
rect 33 -1998 63 -1967
rect -63 -2169 -33 -2138
rect 33 -2164 63 -2138
rect -81 -2185 -15 -2169
rect -81 -2219 -65 -2185
rect -31 -2219 -15 -2185
rect -81 -2235 -15 -2219
rect -81 -2293 -15 -2277
rect -81 -2327 -65 -2293
rect -31 -2327 -15 -2293
rect -81 -2343 -15 -2327
rect -63 -2374 -33 -2343
rect 33 -2374 63 -2348
rect -63 -2540 -33 -2514
rect 33 -2545 63 -2514
rect 15 -2561 81 -2545
rect 15 -2595 31 -2561
rect 65 -2595 81 -2561
rect 15 -2611 81 -2595
rect 15 -2669 81 -2653
rect 15 -2703 31 -2669
rect 65 -2703 81 -2669
rect 15 -2719 81 -2703
rect -63 -2750 -33 -2724
rect 33 -2750 63 -2719
rect -63 -2921 -33 -2890
rect 33 -2916 63 -2890
rect -81 -2937 -15 -2921
rect -81 -2971 -65 -2937
rect -31 -2971 -15 -2937
rect -81 -2987 -15 -2971
<< polycont >>
rect -65 2937 -31 2971
rect 31 2669 65 2703
rect 31 2561 65 2595
rect -65 2293 -31 2327
rect -65 2185 -31 2219
rect 31 1917 65 1951
rect 31 1809 65 1843
rect -65 1541 -31 1575
rect -65 1433 -31 1467
rect 31 1165 65 1199
rect 31 1057 65 1091
rect -65 789 -31 823
rect -65 681 -31 715
rect 31 413 65 447
rect 31 305 65 339
rect -65 37 -31 71
rect -65 -71 -31 -37
rect 31 -339 65 -305
rect 31 -447 65 -413
rect -65 -715 -31 -681
rect -65 -823 -31 -789
rect 31 -1091 65 -1057
rect 31 -1199 65 -1165
rect -65 -1467 -31 -1433
rect -65 -1575 -31 -1541
rect 31 -1843 65 -1809
rect 31 -1951 65 -1917
rect -65 -2219 -31 -2185
rect -65 -2327 -31 -2293
rect 31 -2595 65 -2561
rect 31 -2703 65 -2669
rect -65 -2971 -31 -2937
<< locali >>
rect -227 3039 -131 3073
rect 131 3039 227 3073
rect -227 2977 -193 3039
rect 193 2977 227 3039
rect -81 2937 -65 2971
rect -31 2937 -15 2971
rect -113 2878 -79 2894
rect -113 2746 -79 2762
rect -17 2878 17 2894
rect -17 2746 17 2762
rect 79 2878 113 2894
rect 79 2746 113 2762
rect 15 2669 31 2703
rect 65 2669 81 2703
rect 15 2561 31 2595
rect 65 2561 81 2595
rect -113 2502 -79 2518
rect -113 2370 -79 2386
rect -17 2502 17 2518
rect -17 2370 17 2386
rect 79 2502 113 2518
rect 79 2370 113 2386
rect -81 2293 -65 2327
rect -31 2293 -15 2327
rect -81 2185 -65 2219
rect -31 2185 -15 2219
rect -113 2126 -79 2142
rect -113 1994 -79 2010
rect -17 2126 17 2142
rect -17 1994 17 2010
rect 79 2126 113 2142
rect 79 1994 113 2010
rect 15 1917 31 1951
rect 65 1917 81 1951
rect 15 1809 31 1843
rect 65 1809 81 1843
rect -113 1750 -79 1766
rect -113 1618 -79 1634
rect -17 1750 17 1766
rect -17 1618 17 1634
rect 79 1750 113 1766
rect 79 1618 113 1634
rect -81 1541 -65 1575
rect -31 1541 -15 1575
rect -81 1433 -65 1467
rect -31 1433 -15 1467
rect -113 1374 -79 1390
rect -113 1242 -79 1258
rect -17 1374 17 1390
rect -17 1242 17 1258
rect 79 1374 113 1390
rect 79 1242 113 1258
rect 15 1165 31 1199
rect 65 1165 81 1199
rect 15 1057 31 1091
rect 65 1057 81 1091
rect -113 998 -79 1014
rect -113 866 -79 882
rect -17 998 17 1014
rect -17 866 17 882
rect 79 998 113 1014
rect 79 866 113 882
rect -81 789 -65 823
rect -31 789 -15 823
rect -81 681 -65 715
rect -31 681 -15 715
rect -113 622 -79 638
rect -113 490 -79 506
rect -17 622 17 638
rect -17 490 17 506
rect 79 622 113 638
rect 79 490 113 506
rect 15 413 31 447
rect 65 413 81 447
rect 15 305 31 339
rect 65 305 81 339
rect -113 246 -79 262
rect -113 114 -79 130
rect -17 246 17 262
rect -17 114 17 130
rect 79 246 113 262
rect 79 114 113 130
rect -81 37 -65 71
rect -31 37 -15 71
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect -113 -130 -79 -114
rect -113 -262 -79 -246
rect -17 -130 17 -114
rect -17 -262 17 -246
rect 79 -130 113 -114
rect 79 -262 113 -246
rect 15 -339 31 -305
rect 65 -339 81 -305
rect 15 -447 31 -413
rect 65 -447 81 -413
rect -113 -506 -79 -490
rect -113 -638 -79 -622
rect -17 -506 17 -490
rect -17 -638 17 -622
rect 79 -506 113 -490
rect 79 -638 113 -622
rect -81 -715 -65 -681
rect -31 -715 -15 -681
rect -81 -823 -65 -789
rect -31 -823 -15 -789
rect -113 -882 -79 -866
rect -113 -1014 -79 -998
rect -17 -882 17 -866
rect -17 -1014 17 -998
rect 79 -882 113 -866
rect 79 -1014 113 -998
rect 15 -1091 31 -1057
rect 65 -1091 81 -1057
rect 15 -1199 31 -1165
rect 65 -1199 81 -1165
rect -113 -1258 -79 -1242
rect -113 -1390 -79 -1374
rect -17 -1258 17 -1242
rect -17 -1390 17 -1374
rect 79 -1258 113 -1242
rect 79 -1390 113 -1374
rect -81 -1467 -65 -1433
rect -31 -1467 -15 -1433
rect -81 -1575 -65 -1541
rect -31 -1575 -15 -1541
rect -113 -1634 -79 -1618
rect -113 -1766 -79 -1750
rect -17 -1634 17 -1618
rect -17 -1766 17 -1750
rect 79 -1634 113 -1618
rect 79 -1766 113 -1750
rect 15 -1843 31 -1809
rect 65 -1843 81 -1809
rect 15 -1951 31 -1917
rect 65 -1951 81 -1917
rect -113 -2010 -79 -1994
rect -113 -2142 -79 -2126
rect -17 -2010 17 -1994
rect -17 -2142 17 -2126
rect 79 -2010 113 -1994
rect 79 -2142 113 -2126
rect -81 -2219 -65 -2185
rect -31 -2219 -15 -2185
rect -81 -2327 -65 -2293
rect -31 -2327 -15 -2293
rect -113 -2386 -79 -2370
rect -113 -2518 -79 -2502
rect -17 -2386 17 -2370
rect -17 -2518 17 -2502
rect 79 -2386 113 -2370
rect 79 -2518 113 -2502
rect 15 -2595 31 -2561
rect 65 -2595 81 -2561
rect 15 -2703 31 -2669
rect 65 -2703 81 -2669
rect -113 -2762 -79 -2746
rect -113 -2894 -79 -2878
rect -17 -2762 17 -2746
rect -17 -2894 17 -2878
rect 79 -2762 113 -2746
rect 79 -2894 113 -2878
rect -81 -2971 -65 -2937
rect -31 -2971 -15 -2937
rect -227 -3039 -193 -2977
rect 193 -3039 227 -2977
rect -227 -3073 -131 -3039
rect 131 -3073 227 -3039
<< viali >>
rect -65 2937 -31 2971
rect -113 2762 -79 2878
rect -17 2762 17 2878
rect 79 2762 113 2878
rect 31 2669 65 2703
rect 31 2561 65 2595
rect -113 2386 -79 2502
rect -17 2386 17 2502
rect 79 2386 113 2502
rect -65 2293 -31 2327
rect -65 2185 -31 2219
rect -113 2010 -79 2126
rect -17 2010 17 2126
rect 79 2010 113 2126
rect 31 1917 65 1951
rect 31 1809 65 1843
rect -113 1634 -79 1750
rect -17 1634 17 1750
rect 79 1634 113 1750
rect -65 1541 -31 1575
rect -65 1433 -31 1467
rect -113 1258 -79 1374
rect -17 1258 17 1374
rect 79 1258 113 1374
rect 31 1165 65 1199
rect 31 1057 65 1091
rect -113 882 -79 998
rect -17 882 17 998
rect 79 882 113 998
rect -65 789 -31 823
rect -65 681 -31 715
rect -113 506 -79 622
rect -17 506 17 622
rect 79 506 113 622
rect 31 413 65 447
rect 31 305 65 339
rect -113 130 -79 246
rect -17 130 17 246
rect 79 130 113 246
rect -65 37 -31 71
rect -65 -71 -31 -37
rect -113 -246 -79 -130
rect -17 -246 17 -130
rect 79 -246 113 -130
rect 31 -339 65 -305
rect 31 -447 65 -413
rect -113 -622 -79 -506
rect -17 -622 17 -506
rect 79 -622 113 -506
rect -65 -715 -31 -681
rect -65 -823 -31 -789
rect -113 -998 -79 -882
rect -17 -998 17 -882
rect 79 -998 113 -882
rect 31 -1091 65 -1057
rect 31 -1199 65 -1165
rect -113 -1374 -79 -1258
rect -17 -1374 17 -1258
rect 79 -1374 113 -1258
rect -65 -1467 -31 -1433
rect -65 -1575 -31 -1541
rect -113 -1750 -79 -1634
rect -17 -1750 17 -1634
rect 79 -1750 113 -1634
rect 31 -1843 65 -1809
rect 31 -1951 65 -1917
rect -113 -2126 -79 -2010
rect -17 -2126 17 -2010
rect 79 -2126 113 -2010
rect -65 -2219 -31 -2185
rect -65 -2327 -31 -2293
rect -113 -2502 -79 -2386
rect -17 -2502 17 -2386
rect 79 -2502 113 -2386
rect 31 -2595 65 -2561
rect 31 -2703 65 -2669
rect -113 -2878 -79 -2762
rect -17 -2878 17 -2762
rect 79 -2878 113 -2762
rect -65 -2971 -31 -2937
<< metal1 >>
rect -77 2971 -19 2977
rect -77 2937 -65 2971
rect -31 2937 -19 2971
rect -77 2931 -19 2937
rect -119 2878 -73 2890
rect -119 2762 -113 2878
rect -79 2762 -73 2878
rect -119 2750 -73 2762
rect -23 2878 23 2890
rect -23 2762 -17 2878
rect 17 2762 23 2878
rect -23 2750 23 2762
rect 73 2878 119 2890
rect 73 2762 79 2878
rect 113 2762 119 2878
rect 73 2750 119 2762
rect 19 2703 77 2709
rect 19 2669 31 2703
rect 65 2669 77 2703
rect 19 2663 77 2669
rect 19 2595 77 2601
rect 19 2561 31 2595
rect 65 2561 77 2595
rect 19 2555 77 2561
rect -119 2502 -73 2514
rect -119 2386 -113 2502
rect -79 2386 -73 2502
rect -119 2374 -73 2386
rect -23 2502 23 2514
rect -23 2386 -17 2502
rect 17 2386 23 2502
rect -23 2374 23 2386
rect 73 2502 119 2514
rect 73 2386 79 2502
rect 113 2386 119 2502
rect 73 2374 119 2386
rect -77 2327 -19 2333
rect -77 2293 -65 2327
rect -31 2293 -19 2327
rect -77 2287 -19 2293
rect -77 2219 -19 2225
rect -77 2185 -65 2219
rect -31 2185 -19 2219
rect -77 2179 -19 2185
rect -119 2126 -73 2138
rect -119 2010 -113 2126
rect -79 2010 -73 2126
rect -119 1998 -73 2010
rect -23 2126 23 2138
rect -23 2010 -17 2126
rect 17 2010 23 2126
rect -23 1998 23 2010
rect 73 2126 119 2138
rect 73 2010 79 2126
rect 113 2010 119 2126
rect 73 1998 119 2010
rect 19 1951 77 1957
rect 19 1917 31 1951
rect 65 1917 77 1951
rect 19 1911 77 1917
rect 19 1843 77 1849
rect 19 1809 31 1843
rect 65 1809 77 1843
rect 19 1803 77 1809
rect -119 1750 -73 1762
rect -119 1634 -113 1750
rect -79 1634 -73 1750
rect -119 1622 -73 1634
rect -23 1750 23 1762
rect -23 1634 -17 1750
rect 17 1634 23 1750
rect -23 1622 23 1634
rect 73 1750 119 1762
rect 73 1634 79 1750
rect 113 1634 119 1750
rect 73 1622 119 1634
rect -77 1575 -19 1581
rect -77 1541 -65 1575
rect -31 1541 -19 1575
rect -77 1535 -19 1541
rect -77 1467 -19 1473
rect -77 1433 -65 1467
rect -31 1433 -19 1467
rect -77 1427 -19 1433
rect -119 1374 -73 1386
rect -119 1258 -113 1374
rect -79 1258 -73 1374
rect -119 1246 -73 1258
rect -23 1374 23 1386
rect -23 1258 -17 1374
rect 17 1258 23 1374
rect -23 1246 23 1258
rect 73 1374 119 1386
rect 73 1258 79 1374
rect 113 1258 119 1374
rect 73 1246 119 1258
rect 19 1199 77 1205
rect 19 1165 31 1199
rect 65 1165 77 1199
rect 19 1159 77 1165
rect 19 1091 77 1097
rect 19 1057 31 1091
rect 65 1057 77 1091
rect 19 1051 77 1057
rect -119 998 -73 1010
rect -119 882 -113 998
rect -79 882 -73 998
rect -119 870 -73 882
rect -23 998 23 1010
rect -23 882 -17 998
rect 17 882 23 998
rect -23 870 23 882
rect 73 998 119 1010
rect 73 882 79 998
rect 113 882 119 998
rect 73 870 119 882
rect -77 823 -19 829
rect -77 789 -65 823
rect -31 789 -19 823
rect -77 783 -19 789
rect -77 715 -19 721
rect -77 681 -65 715
rect -31 681 -19 715
rect -77 675 -19 681
rect -119 622 -73 634
rect -119 506 -113 622
rect -79 506 -73 622
rect -119 494 -73 506
rect -23 622 23 634
rect -23 506 -17 622
rect 17 506 23 622
rect -23 494 23 506
rect 73 622 119 634
rect 73 506 79 622
rect 113 506 119 622
rect 73 494 119 506
rect 19 447 77 453
rect 19 413 31 447
rect 65 413 77 447
rect 19 407 77 413
rect 19 339 77 345
rect 19 305 31 339
rect 65 305 77 339
rect 19 299 77 305
rect -119 246 -73 258
rect -119 130 -113 246
rect -79 130 -73 246
rect -119 118 -73 130
rect -23 246 23 258
rect -23 130 -17 246
rect 17 130 23 246
rect -23 118 23 130
rect 73 246 119 258
rect 73 130 79 246
rect 113 130 119 246
rect 73 118 119 130
rect -77 71 -19 77
rect -77 37 -65 71
rect -31 37 -19 71
rect -77 31 -19 37
rect -77 -37 -19 -31
rect -77 -71 -65 -37
rect -31 -71 -19 -37
rect -77 -77 -19 -71
rect -119 -130 -73 -118
rect -119 -246 -113 -130
rect -79 -246 -73 -130
rect -119 -258 -73 -246
rect -23 -130 23 -118
rect -23 -246 -17 -130
rect 17 -246 23 -130
rect -23 -258 23 -246
rect 73 -130 119 -118
rect 73 -246 79 -130
rect 113 -246 119 -130
rect 73 -258 119 -246
rect 19 -305 77 -299
rect 19 -339 31 -305
rect 65 -339 77 -305
rect 19 -345 77 -339
rect 19 -413 77 -407
rect 19 -447 31 -413
rect 65 -447 77 -413
rect 19 -453 77 -447
rect -119 -506 -73 -494
rect -119 -622 -113 -506
rect -79 -622 -73 -506
rect -119 -634 -73 -622
rect -23 -506 23 -494
rect -23 -622 -17 -506
rect 17 -622 23 -506
rect -23 -634 23 -622
rect 73 -506 119 -494
rect 73 -622 79 -506
rect 113 -622 119 -506
rect 73 -634 119 -622
rect -77 -681 -19 -675
rect -77 -715 -65 -681
rect -31 -715 -19 -681
rect -77 -721 -19 -715
rect -77 -789 -19 -783
rect -77 -823 -65 -789
rect -31 -823 -19 -789
rect -77 -829 -19 -823
rect -119 -882 -73 -870
rect -119 -998 -113 -882
rect -79 -998 -73 -882
rect -119 -1010 -73 -998
rect -23 -882 23 -870
rect -23 -998 -17 -882
rect 17 -998 23 -882
rect -23 -1010 23 -998
rect 73 -882 119 -870
rect 73 -998 79 -882
rect 113 -998 119 -882
rect 73 -1010 119 -998
rect 19 -1057 77 -1051
rect 19 -1091 31 -1057
rect 65 -1091 77 -1057
rect 19 -1097 77 -1091
rect 19 -1165 77 -1159
rect 19 -1199 31 -1165
rect 65 -1199 77 -1165
rect 19 -1205 77 -1199
rect -119 -1258 -73 -1246
rect -119 -1374 -113 -1258
rect -79 -1374 -73 -1258
rect -119 -1386 -73 -1374
rect -23 -1258 23 -1246
rect -23 -1374 -17 -1258
rect 17 -1374 23 -1258
rect -23 -1386 23 -1374
rect 73 -1258 119 -1246
rect 73 -1374 79 -1258
rect 113 -1374 119 -1258
rect 73 -1386 119 -1374
rect -77 -1433 -19 -1427
rect -77 -1467 -65 -1433
rect -31 -1467 -19 -1433
rect -77 -1473 -19 -1467
rect -77 -1541 -19 -1535
rect -77 -1575 -65 -1541
rect -31 -1575 -19 -1541
rect -77 -1581 -19 -1575
rect -119 -1634 -73 -1622
rect -119 -1750 -113 -1634
rect -79 -1750 -73 -1634
rect -119 -1762 -73 -1750
rect -23 -1634 23 -1622
rect -23 -1750 -17 -1634
rect 17 -1750 23 -1634
rect -23 -1762 23 -1750
rect 73 -1634 119 -1622
rect 73 -1750 79 -1634
rect 113 -1750 119 -1634
rect 73 -1762 119 -1750
rect 19 -1809 77 -1803
rect 19 -1843 31 -1809
rect 65 -1843 77 -1809
rect 19 -1849 77 -1843
rect 19 -1917 77 -1911
rect 19 -1951 31 -1917
rect 65 -1951 77 -1917
rect 19 -1957 77 -1951
rect -119 -2010 -73 -1998
rect -119 -2126 -113 -2010
rect -79 -2126 -73 -2010
rect -119 -2138 -73 -2126
rect -23 -2010 23 -1998
rect -23 -2126 -17 -2010
rect 17 -2126 23 -2010
rect -23 -2138 23 -2126
rect 73 -2010 119 -1998
rect 73 -2126 79 -2010
rect 113 -2126 119 -2010
rect 73 -2138 119 -2126
rect -77 -2185 -19 -2179
rect -77 -2219 -65 -2185
rect -31 -2219 -19 -2185
rect -77 -2225 -19 -2219
rect -77 -2293 -19 -2287
rect -77 -2327 -65 -2293
rect -31 -2327 -19 -2293
rect -77 -2333 -19 -2327
rect -119 -2386 -73 -2374
rect -119 -2502 -113 -2386
rect -79 -2502 -73 -2386
rect -119 -2514 -73 -2502
rect -23 -2386 23 -2374
rect -23 -2502 -17 -2386
rect 17 -2502 23 -2386
rect -23 -2514 23 -2502
rect 73 -2386 119 -2374
rect 73 -2502 79 -2386
rect 113 -2502 119 -2386
rect 73 -2514 119 -2502
rect 19 -2561 77 -2555
rect 19 -2595 31 -2561
rect 65 -2595 77 -2561
rect 19 -2601 77 -2595
rect 19 -2669 77 -2663
rect 19 -2703 31 -2669
rect 65 -2703 77 -2669
rect 19 -2709 77 -2703
rect -119 -2762 -73 -2750
rect -119 -2878 -113 -2762
rect -79 -2878 -73 -2762
rect -119 -2890 -73 -2878
rect -23 -2762 23 -2750
rect -23 -2878 -17 -2762
rect 17 -2878 23 -2762
rect -23 -2890 23 -2878
rect 73 -2762 119 -2750
rect 73 -2878 79 -2762
rect 113 -2878 119 -2762
rect 73 -2890 119 -2878
rect -77 -2937 -19 -2931
rect -77 -2971 -65 -2937
rect -31 -2971 -19 -2937
rect -77 -2977 -19 -2971
<< properties >>
string FIXED_BBOX -210 -3056 210 3056
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.7 l 0.15 m 16 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
