magic
tech sky130A
magscale 1 2
timestamp 1717363523
<< metal4 >>
rect -8396 17839 -4498 17880
rect -8396 14561 -4754 17839
rect -4518 14561 -4498 17839
rect -8396 14520 -4498 14561
rect -4098 17839 -200 17880
rect -4098 14561 -456 17839
rect -220 14561 -200 17839
rect -4098 14520 -200 14561
rect 200 17839 4098 17880
rect 200 14561 3842 17839
rect 4078 14561 4098 17839
rect 200 14520 4098 14561
rect 4498 17839 8396 17880
rect 4498 14561 8140 17839
rect 8376 14561 8396 17839
rect 4498 14520 8396 14561
rect -8396 14239 -4498 14280
rect -8396 10961 -4754 14239
rect -4518 10961 -4498 14239
rect -8396 10920 -4498 10961
rect -4098 14239 -200 14280
rect -4098 10961 -456 14239
rect -220 10961 -200 14239
rect -4098 10920 -200 10961
rect 200 14239 4098 14280
rect 200 10961 3842 14239
rect 4078 10961 4098 14239
rect 200 10920 4098 10961
rect 4498 14239 8396 14280
rect 4498 10961 8140 14239
rect 8376 10961 8396 14239
rect 4498 10920 8396 10961
rect -8396 10639 -4498 10680
rect -8396 7361 -4754 10639
rect -4518 7361 -4498 10639
rect -8396 7320 -4498 7361
rect -4098 10639 -200 10680
rect -4098 7361 -456 10639
rect -220 7361 -200 10639
rect -4098 7320 -200 7361
rect 200 10639 4098 10680
rect 200 7361 3842 10639
rect 4078 7361 4098 10639
rect 200 7320 4098 7361
rect 4498 10639 8396 10680
rect 4498 7361 8140 10639
rect 8376 7361 8396 10639
rect 4498 7320 8396 7361
rect -8396 7039 -4498 7080
rect -8396 3761 -4754 7039
rect -4518 3761 -4498 7039
rect -8396 3720 -4498 3761
rect -4098 7039 -200 7080
rect -4098 3761 -456 7039
rect -220 3761 -200 7039
rect -4098 3720 -200 3761
rect 200 7039 4098 7080
rect 200 3761 3842 7039
rect 4078 3761 4098 7039
rect 200 3720 4098 3761
rect 4498 7039 8396 7080
rect 4498 3761 8140 7039
rect 8376 3761 8396 7039
rect 4498 3720 8396 3761
rect -8396 3439 -4498 3480
rect -8396 161 -4754 3439
rect -4518 161 -4498 3439
rect -8396 120 -4498 161
rect -4098 3439 -200 3480
rect -4098 161 -456 3439
rect -220 161 -200 3439
rect -4098 120 -200 161
rect 200 3439 4098 3480
rect 200 161 3842 3439
rect 4078 161 4098 3439
rect 200 120 4098 161
rect 4498 3439 8396 3480
rect 4498 161 8140 3439
rect 8376 161 8396 3439
rect 4498 120 8396 161
rect -8396 -161 -4498 -120
rect -8396 -3439 -4754 -161
rect -4518 -3439 -4498 -161
rect -8396 -3480 -4498 -3439
rect -4098 -161 -200 -120
rect -4098 -3439 -456 -161
rect -220 -3439 -200 -161
rect -4098 -3480 -200 -3439
rect 200 -161 4098 -120
rect 200 -3439 3842 -161
rect 4078 -3439 4098 -161
rect 200 -3480 4098 -3439
rect 4498 -161 8396 -120
rect 4498 -3439 8140 -161
rect 8376 -3439 8396 -161
rect 4498 -3480 8396 -3439
rect -8396 -3761 -4498 -3720
rect -8396 -7039 -4754 -3761
rect -4518 -7039 -4498 -3761
rect -8396 -7080 -4498 -7039
rect -4098 -3761 -200 -3720
rect -4098 -7039 -456 -3761
rect -220 -7039 -200 -3761
rect -4098 -7080 -200 -7039
rect 200 -3761 4098 -3720
rect 200 -7039 3842 -3761
rect 4078 -7039 4098 -3761
rect 200 -7080 4098 -7039
rect 4498 -3761 8396 -3720
rect 4498 -7039 8140 -3761
rect 8376 -7039 8396 -3761
rect 4498 -7080 8396 -7039
rect -8396 -7361 -4498 -7320
rect -8396 -10639 -4754 -7361
rect -4518 -10639 -4498 -7361
rect -8396 -10680 -4498 -10639
rect -4098 -7361 -200 -7320
rect -4098 -10639 -456 -7361
rect -220 -10639 -200 -7361
rect -4098 -10680 -200 -10639
rect 200 -7361 4098 -7320
rect 200 -10639 3842 -7361
rect 4078 -10639 4098 -7361
rect 200 -10680 4098 -10639
rect 4498 -7361 8396 -7320
rect 4498 -10639 8140 -7361
rect 8376 -10639 8396 -7361
rect 4498 -10680 8396 -10639
rect -8396 -10961 -4498 -10920
rect -8396 -14239 -4754 -10961
rect -4518 -14239 -4498 -10961
rect -8396 -14280 -4498 -14239
rect -4098 -10961 -200 -10920
rect -4098 -14239 -456 -10961
rect -220 -14239 -200 -10961
rect -4098 -14280 -200 -14239
rect 200 -10961 4098 -10920
rect 200 -14239 3842 -10961
rect 4078 -14239 4098 -10961
rect 200 -14280 4098 -14239
rect 4498 -10961 8396 -10920
rect 4498 -14239 8140 -10961
rect 8376 -14239 8396 -10961
rect 4498 -14280 8396 -14239
rect -8396 -14561 -4498 -14520
rect -8396 -17839 -4754 -14561
rect -4518 -17839 -4498 -14561
rect -8396 -17880 -4498 -17839
rect -4098 -14561 -200 -14520
rect -4098 -17839 -456 -14561
rect -220 -17839 -200 -14561
rect -4098 -17880 -200 -17839
rect 200 -14561 4098 -14520
rect 200 -17839 3842 -14561
rect 4078 -17839 4098 -14561
rect 200 -17880 4098 -17839
rect 4498 -14561 8396 -14520
rect 4498 -17839 8140 -14561
rect 8376 -17839 8396 -14561
rect 4498 -17880 8396 -17839
<< via4 >>
rect -4754 14561 -4518 17839
rect -456 14561 -220 17839
rect 3842 14561 4078 17839
rect 8140 14561 8376 17839
rect -4754 10961 -4518 14239
rect -456 10961 -220 14239
rect 3842 10961 4078 14239
rect 8140 10961 8376 14239
rect -4754 7361 -4518 10639
rect -456 7361 -220 10639
rect 3842 7361 4078 10639
rect 8140 7361 8376 10639
rect -4754 3761 -4518 7039
rect -456 3761 -220 7039
rect 3842 3761 4078 7039
rect 8140 3761 8376 7039
rect -4754 161 -4518 3439
rect -456 161 -220 3439
rect 3842 161 4078 3439
rect 8140 161 8376 3439
rect -4754 -3439 -4518 -161
rect -456 -3439 -220 -161
rect 3842 -3439 4078 -161
rect 8140 -3439 8376 -161
rect -4754 -7039 -4518 -3761
rect -456 -7039 -220 -3761
rect 3842 -7039 4078 -3761
rect 8140 -7039 8376 -3761
rect -4754 -10639 -4518 -7361
rect -456 -10639 -220 -7361
rect 3842 -10639 4078 -7361
rect 8140 -10639 8376 -7361
rect -4754 -14239 -4518 -10961
rect -456 -14239 -220 -10961
rect 3842 -14239 4078 -10961
rect 8140 -14239 8376 -10961
rect -4754 -17839 -4518 -14561
rect -456 -17839 -220 -14561
rect 3842 -17839 4078 -14561
rect 8140 -17839 8376 -14561
<< mimcap2 >>
rect -8316 17760 -5116 17800
rect -8316 14640 -8276 17760
rect -5156 14640 -5116 17760
rect -8316 14600 -5116 14640
rect -4018 17760 -818 17800
rect -4018 14640 -3978 17760
rect -858 14640 -818 17760
rect -4018 14600 -818 14640
rect 280 17760 3480 17800
rect 280 14640 320 17760
rect 3440 14640 3480 17760
rect 280 14600 3480 14640
rect 4578 17760 7778 17800
rect 4578 14640 4618 17760
rect 7738 14640 7778 17760
rect 4578 14600 7778 14640
rect -8316 14160 -5116 14200
rect -8316 11040 -8276 14160
rect -5156 11040 -5116 14160
rect -8316 11000 -5116 11040
rect -4018 14160 -818 14200
rect -4018 11040 -3978 14160
rect -858 11040 -818 14160
rect -4018 11000 -818 11040
rect 280 14160 3480 14200
rect 280 11040 320 14160
rect 3440 11040 3480 14160
rect 280 11000 3480 11040
rect 4578 14160 7778 14200
rect 4578 11040 4618 14160
rect 7738 11040 7778 14160
rect 4578 11000 7778 11040
rect -8316 10560 -5116 10600
rect -8316 7440 -8276 10560
rect -5156 7440 -5116 10560
rect -8316 7400 -5116 7440
rect -4018 10560 -818 10600
rect -4018 7440 -3978 10560
rect -858 7440 -818 10560
rect -4018 7400 -818 7440
rect 280 10560 3480 10600
rect 280 7440 320 10560
rect 3440 7440 3480 10560
rect 280 7400 3480 7440
rect 4578 10560 7778 10600
rect 4578 7440 4618 10560
rect 7738 7440 7778 10560
rect 4578 7400 7778 7440
rect -8316 6960 -5116 7000
rect -8316 3840 -8276 6960
rect -5156 3840 -5116 6960
rect -8316 3800 -5116 3840
rect -4018 6960 -818 7000
rect -4018 3840 -3978 6960
rect -858 3840 -818 6960
rect -4018 3800 -818 3840
rect 280 6960 3480 7000
rect 280 3840 320 6960
rect 3440 3840 3480 6960
rect 280 3800 3480 3840
rect 4578 6960 7778 7000
rect 4578 3840 4618 6960
rect 7738 3840 7778 6960
rect 4578 3800 7778 3840
rect -8316 3360 -5116 3400
rect -8316 240 -8276 3360
rect -5156 240 -5116 3360
rect -8316 200 -5116 240
rect -4018 3360 -818 3400
rect -4018 240 -3978 3360
rect -858 240 -818 3360
rect -4018 200 -818 240
rect 280 3360 3480 3400
rect 280 240 320 3360
rect 3440 240 3480 3360
rect 280 200 3480 240
rect 4578 3360 7778 3400
rect 4578 240 4618 3360
rect 7738 240 7778 3360
rect 4578 200 7778 240
rect -8316 -240 -5116 -200
rect -8316 -3360 -8276 -240
rect -5156 -3360 -5116 -240
rect -8316 -3400 -5116 -3360
rect -4018 -240 -818 -200
rect -4018 -3360 -3978 -240
rect -858 -3360 -818 -240
rect -4018 -3400 -818 -3360
rect 280 -240 3480 -200
rect 280 -3360 320 -240
rect 3440 -3360 3480 -240
rect 280 -3400 3480 -3360
rect 4578 -240 7778 -200
rect 4578 -3360 4618 -240
rect 7738 -3360 7778 -240
rect 4578 -3400 7778 -3360
rect -8316 -3840 -5116 -3800
rect -8316 -6960 -8276 -3840
rect -5156 -6960 -5116 -3840
rect -8316 -7000 -5116 -6960
rect -4018 -3840 -818 -3800
rect -4018 -6960 -3978 -3840
rect -858 -6960 -818 -3840
rect -4018 -7000 -818 -6960
rect 280 -3840 3480 -3800
rect 280 -6960 320 -3840
rect 3440 -6960 3480 -3840
rect 280 -7000 3480 -6960
rect 4578 -3840 7778 -3800
rect 4578 -6960 4618 -3840
rect 7738 -6960 7778 -3840
rect 4578 -7000 7778 -6960
rect -8316 -7440 -5116 -7400
rect -8316 -10560 -8276 -7440
rect -5156 -10560 -5116 -7440
rect -8316 -10600 -5116 -10560
rect -4018 -7440 -818 -7400
rect -4018 -10560 -3978 -7440
rect -858 -10560 -818 -7440
rect -4018 -10600 -818 -10560
rect 280 -7440 3480 -7400
rect 280 -10560 320 -7440
rect 3440 -10560 3480 -7440
rect 280 -10600 3480 -10560
rect 4578 -7440 7778 -7400
rect 4578 -10560 4618 -7440
rect 7738 -10560 7778 -7440
rect 4578 -10600 7778 -10560
rect -8316 -11040 -5116 -11000
rect -8316 -14160 -8276 -11040
rect -5156 -14160 -5116 -11040
rect -8316 -14200 -5116 -14160
rect -4018 -11040 -818 -11000
rect -4018 -14160 -3978 -11040
rect -858 -14160 -818 -11040
rect -4018 -14200 -818 -14160
rect 280 -11040 3480 -11000
rect 280 -14160 320 -11040
rect 3440 -14160 3480 -11040
rect 280 -14200 3480 -14160
rect 4578 -11040 7778 -11000
rect 4578 -14160 4618 -11040
rect 7738 -14160 7778 -11040
rect 4578 -14200 7778 -14160
rect -8316 -14640 -5116 -14600
rect -8316 -17760 -8276 -14640
rect -5156 -17760 -5116 -14640
rect -8316 -17800 -5116 -17760
rect -4018 -14640 -818 -14600
rect -4018 -17760 -3978 -14640
rect -858 -17760 -818 -14640
rect -4018 -17800 -818 -17760
rect 280 -14640 3480 -14600
rect 280 -17760 320 -14640
rect 3440 -17760 3480 -14640
rect 280 -17800 3480 -17760
rect 4578 -14640 7778 -14600
rect 4578 -17760 4618 -14640
rect 7738 -17760 7778 -14640
rect 4578 -17800 7778 -17760
<< mimcap2contact >>
rect -8276 14640 -5156 17760
rect -3978 14640 -858 17760
rect 320 14640 3440 17760
rect 4618 14640 7738 17760
rect -8276 11040 -5156 14160
rect -3978 11040 -858 14160
rect 320 11040 3440 14160
rect 4618 11040 7738 14160
rect -8276 7440 -5156 10560
rect -3978 7440 -858 10560
rect 320 7440 3440 10560
rect 4618 7440 7738 10560
rect -8276 3840 -5156 6960
rect -3978 3840 -858 6960
rect 320 3840 3440 6960
rect 4618 3840 7738 6960
rect -8276 240 -5156 3360
rect -3978 240 -858 3360
rect 320 240 3440 3360
rect 4618 240 7738 3360
rect -8276 -3360 -5156 -240
rect -3978 -3360 -858 -240
rect 320 -3360 3440 -240
rect 4618 -3360 7738 -240
rect -8276 -6960 -5156 -3840
rect -3978 -6960 -858 -3840
rect 320 -6960 3440 -3840
rect 4618 -6960 7738 -3840
rect -8276 -10560 -5156 -7440
rect -3978 -10560 -858 -7440
rect 320 -10560 3440 -7440
rect 4618 -10560 7738 -7440
rect -8276 -14160 -5156 -11040
rect -3978 -14160 -858 -11040
rect 320 -14160 3440 -11040
rect 4618 -14160 7738 -11040
rect -8276 -17760 -5156 -14640
rect -3978 -17760 -858 -14640
rect 320 -17760 3440 -14640
rect 4618 -17760 7738 -14640
<< metal5 >>
rect -6876 17784 -6556 18000
rect -4796 17839 -4476 18000
rect -8300 17760 -5132 17784
rect -8300 14640 -8276 17760
rect -5156 14640 -5132 17760
rect -8300 14616 -5132 14640
rect -6876 14184 -6556 14616
rect -4796 14561 -4754 17839
rect -4518 14561 -4476 17839
rect -2578 17784 -2258 18000
rect -498 17839 -178 18000
rect -4002 17760 -834 17784
rect -4002 14640 -3978 17760
rect -858 14640 -834 17760
rect -4002 14616 -834 14640
rect -4796 14239 -4476 14561
rect -8300 14160 -5132 14184
rect -8300 11040 -8276 14160
rect -5156 11040 -5132 14160
rect -8300 11016 -5132 11040
rect -6876 10584 -6556 11016
rect -4796 10961 -4754 14239
rect -4518 10961 -4476 14239
rect -2578 14184 -2258 14616
rect -498 14561 -456 17839
rect -220 14561 -178 17839
rect 1720 17784 2040 18000
rect 3800 17839 4120 18000
rect 296 17760 3464 17784
rect 296 14640 320 17760
rect 3440 14640 3464 17760
rect 296 14616 3464 14640
rect -498 14239 -178 14561
rect -4002 14160 -834 14184
rect -4002 11040 -3978 14160
rect -858 11040 -834 14160
rect -4002 11016 -834 11040
rect -4796 10639 -4476 10961
rect -8300 10560 -5132 10584
rect -8300 7440 -8276 10560
rect -5156 7440 -5132 10560
rect -8300 7416 -5132 7440
rect -6876 6984 -6556 7416
rect -4796 7361 -4754 10639
rect -4518 7361 -4476 10639
rect -2578 10584 -2258 11016
rect -498 10961 -456 14239
rect -220 10961 -178 14239
rect 1720 14184 2040 14616
rect 3800 14561 3842 17839
rect 4078 14561 4120 17839
rect 6018 17784 6338 18000
rect 8098 17839 8418 18000
rect 4594 17760 7762 17784
rect 4594 14640 4618 17760
rect 7738 14640 7762 17760
rect 4594 14616 7762 14640
rect 3800 14239 4120 14561
rect 296 14160 3464 14184
rect 296 11040 320 14160
rect 3440 11040 3464 14160
rect 296 11016 3464 11040
rect -498 10639 -178 10961
rect -4002 10560 -834 10584
rect -4002 7440 -3978 10560
rect -858 7440 -834 10560
rect -4002 7416 -834 7440
rect -4796 7039 -4476 7361
rect -8300 6960 -5132 6984
rect -8300 3840 -8276 6960
rect -5156 3840 -5132 6960
rect -8300 3816 -5132 3840
rect -6876 3384 -6556 3816
rect -4796 3761 -4754 7039
rect -4518 3761 -4476 7039
rect -2578 6984 -2258 7416
rect -498 7361 -456 10639
rect -220 7361 -178 10639
rect 1720 10584 2040 11016
rect 3800 10961 3842 14239
rect 4078 10961 4120 14239
rect 6018 14184 6338 14616
rect 8098 14561 8140 17839
rect 8376 14561 8418 17839
rect 8098 14239 8418 14561
rect 4594 14160 7762 14184
rect 4594 11040 4618 14160
rect 7738 11040 7762 14160
rect 4594 11016 7762 11040
rect 3800 10639 4120 10961
rect 296 10560 3464 10584
rect 296 7440 320 10560
rect 3440 7440 3464 10560
rect 296 7416 3464 7440
rect -498 7039 -178 7361
rect -4002 6960 -834 6984
rect -4002 3840 -3978 6960
rect -858 3840 -834 6960
rect -4002 3816 -834 3840
rect -4796 3439 -4476 3761
rect -8300 3360 -5132 3384
rect -8300 240 -8276 3360
rect -5156 240 -5132 3360
rect -8300 216 -5132 240
rect -6876 -216 -6556 216
rect -4796 161 -4754 3439
rect -4518 161 -4476 3439
rect -2578 3384 -2258 3816
rect -498 3761 -456 7039
rect -220 3761 -178 7039
rect 1720 6984 2040 7416
rect 3800 7361 3842 10639
rect 4078 7361 4120 10639
rect 6018 10584 6338 11016
rect 8098 10961 8140 14239
rect 8376 10961 8418 14239
rect 8098 10639 8418 10961
rect 4594 10560 7762 10584
rect 4594 7440 4618 10560
rect 7738 7440 7762 10560
rect 4594 7416 7762 7440
rect 3800 7039 4120 7361
rect 296 6960 3464 6984
rect 296 3840 320 6960
rect 3440 3840 3464 6960
rect 296 3816 3464 3840
rect -498 3439 -178 3761
rect -4002 3360 -834 3384
rect -4002 240 -3978 3360
rect -858 240 -834 3360
rect -4002 216 -834 240
rect -4796 -161 -4476 161
rect -8300 -240 -5132 -216
rect -8300 -3360 -8276 -240
rect -5156 -3360 -5132 -240
rect -8300 -3384 -5132 -3360
rect -6876 -3816 -6556 -3384
rect -4796 -3439 -4754 -161
rect -4518 -3439 -4476 -161
rect -2578 -216 -2258 216
rect -498 161 -456 3439
rect -220 161 -178 3439
rect 1720 3384 2040 3816
rect 3800 3761 3842 7039
rect 4078 3761 4120 7039
rect 6018 6984 6338 7416
rect 8098 7361 8140 10639
rect 8376 7361 8418 10639
rect 8098 7039 8418 7361
rect 4594 6960 7762 6984
rect 4594 3840 4618 6960
rect 7738 3840 7762 6960
rect 4594 3816 7762 3840
rect 3800 3439 4120 3761
rect 296 3360 3464 3384
rect 296 240 320 3360
rect 3440 240 3464 3360
rect 296 216 3464 240
rect -498 -161 -178 161
rect -4002 -240 -834 -216
rect -4002 -3360 -3978 -240
rect -858 -3360 -834 -240
rect -4002 -3384 -834 -3360
rect -4796 -3761 -4476 -3439
rect -8300 -3840 -5132 -3816
rect -8300 -6960 -8276 -3840
rect -5156 -6960 -5132 -3840
rect -8300 -6984 -5132 -6960
rect -6876 -7416 -6556 -6984
rect -4796 -7039 -4754 -3761
rect -4518 -7039 -4476 -3761
rect -2578 -3816 -2258 -3384
rect -498 -3439 -456 -161
rect -220 -3439 -178 -161
rect 1720 -216 2040 216
rect 3800 161 3842 3439
rect 4078 161 4120 3439
rect 6018 3384 6338 3816
rect 8098 3761 8140 7039
rect 8376 3761 8418 7039
rect 8098 3439 8418 3761
rect 4594 3360 7762 3384
rect 4594 240 4618 3360
rect 7738 240 7762 3360
rect 4594 216 7762 240
rect 3800 -161 4120 161
rect 296 -240 3464 -216
rect 296 -3360 320 -240
rect 3440 -3360 3464 -240
rect 296 -3384 3464 -3360
rect -498 -3761 -178 -3439
rect -4002 -3840 -834 -3816
rect -4002 -6960 -3978 -3840
rect -858 -6960 -834 -3840
rect -4002 -6984 -834 -6960
rect -4796 -7361 -4476 -7039
rect -8300 -7440 -5132 -7416
rect -8300 -10560 -8276 -7440
rect -5156 -10560 -5132 -7440
rect -8300 -10584 -5132 -10560
rect -6876 -11016 -6556 -10584
rect -4796 -10639 -4754 -7361
rect -4518 -10639 -4476 -7361
rect -2578 -7416 -2258 -6984
rect -498 -7039 -456 -3761
rect -220 -7039 -178 -3761
rect 1720 -3816 2040 -3384
rect 3800 -3439 3842 -161
rect 4078 -3439 4120 -161
rect 6018 -216 6338 216
rect 8098 161 8140 3439
rect 8376 161 8418 3439
rect 8098 -161 8418 161
rect 4594 -240 7762 -216
rect 4594 -3360 4618 -240
rect 7738 -3360 7762 -240
rect 4594 -3384 7762 -3360
rect 3800 -3761 4120 -3439
rect 296 -3840 3464 -3816
rect 296 -6960 320 -3840
rect 3440 -6960 3464 -3840
rect 296 -6984 3464 -6960
rect -498 -7361 -178 -7039
rect -4002 -7440 -834 -7416
rect -4002 -10560 -3978 -7440
rect -858 -10560 -834 -7440
rect -4002 -10584 -834 -10560
rect -4796 -10961 -4476 -10639
rect -8300 -11040 -5132 -11016
rect -8300 -14160 -8276 -11040
rect -5156 -14160 -5132 -11040
rect -8300 -14184 -5132 -14160
rect -6876 -14616 -6556 -14184
rect -4796 -14239 -4754 -10961
rect -4518 -14239 -4476 -10961
rect -2578 -11016 -2258 -10584
rect -498 -10639 -456 -7361
rect -220 -10639 -178 -7361
rect 1720 -7416 2040 -6984
rect 3800 -7039 3842 -3761
rect 4078 -7039 4120 -3761
rect 6018 -3816 6338 -3384
rect 8098 -3439 8140 -161
rect 8376 -3439 8418 -161
rect 8098 -3761 8418 -3439
rect 4594 -3840 7762 -3816
rect 4594 -6960 4618 -3840
rect 7738 -6960 7762 -3840
rect 4594 -6984 7762 -6960
rect 3800 -7361 4120 -7039
rect 296 -7440 3464 -7416
rect 296 -10560 320 -7440
rect 3440 -10560 3464 -7440
rect 296 -10584 3464 -10560
rect -498 -10961 -178 -10639
rect -4002 -11040 -834 -11016
rect -4002 -14160 -3978 -11040
rect -858 -14160 -834 -11040
rect -4002 -14184 -834 -14160
rect -4796 -14561 -4476 -14239
rect -8300 -14640 -5132 -14616
rect -8300 -17760 -8276 -14640
rect -5156 -17760 -5132 -14640
rect -8300 -17784 -5132 -17760
rect -6876 -18000 -6556 -17784
rect -4796 -17839 -4754 -14561
rect -4518 -17839 -4476 -14561
rect -2578 -14616 -2258 -14184
rect -498 -14239 -456 -10961
rect -220 -14239 -178 -10961
rect 1720 -11016 2040 -10584
rect 3800 -10639 3842 -7361
rect 4078 -10639 4120 -7361
rect 6018 -7416 6338 -6984
rect 8098 -7039 8140 -3761
rect 8376 -7039 8418 -3761
rect 8098 -7361 8418 -7039
rect 4594 -7440 7762 -7416
rect 4594 -10560 4618 -7440
rect 7738 -10560 7762 -7440
rect 4594 -10584 7762 -10560
rect 3800 -10961 4120 -10639
rect 296 -11040 3464 -11016
rect 296 -14160 320 -11040
rect 3440 -14160 3464 -11040
rect 296 -14184 3464 -14160
rect -498 -14561 -178 -14239
rect -4002 -14640 -834 -14616
rect -4002 -17760 -3978 -14640
rect -858 -17760 -834 -14640
rect -4002 -17784 -834 -17760
rect -4796 -18000 -4476 -17839
rect -2578 -18000 -2258 -17784
rect -498 -17839 -456 -14561
rect -220 -17839 -178 -14561
rect 1720 -14616 2040 -14184
rect 3800 -14239 3842 -10961
rect 4078 -14239 4120 -10961
rect 6018 -11016 6338 -10584
rect 8098 -10639 8140 -7361
rect 8376 -10639 8418 -7361
rect 8098 -10961 8418 -10639
rect 4594 -11040 7762 -11016
rect 4594 -14160 4618 -11040
rect 7738 -14160 7762 -11040
rect 4594 -14184 7762 -14160
rect 3800 -14561 4120 -14239
rect 296 -14640 3464 -14616
rect 296 -17760 320 -14640
rect 3440 -17760 3464 -14640
rect 296 -17784 3464 -17760
rect -498 -18000 -178 -17839
rect 1720 -18000 2040 -17784
rect 3800 -17839 3842 -14561
rect 4078 -17839 4120 -14561
rect 6018 -14616 6338 -14184
rect 8098 -14239 8140 -10961
rect 8376 -14239 8418 -10961
rect 8098 -14561 8418 -14239
rect 4594 -14640 7762 -14616
rect 4594 -17760 4618 -14640
rect 7738 -17760 7762 -14640
rect 4594 -17784 7762 -17760
rect 3800 -18000 4120 -17839
rect 6018 -18000 6338 -17784
rect 8098 -17839 8140 -14561
rect 8376 -17839 8418 -14561
rect 8098 -18000 8418 -17839
<< properties >>
string FIXED_BBOX 4498 14520 7858 17880
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 16.0 l 16.0 val 524.159 carea 2.00 cperi 0.19 nx 4 ny 10 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
