magic
tech sky130A
magscale 1 2
timestamp 1718283729
<< pwell >>
rect -635 -458 635 458
<< mvnmos >>
rect -407 -200 -247 200
rect -189 -200 -29 200
rect 29 -200 189 200
rect 247 -200 407 200
<< mvndiff >>
rect -465 188 -407 200
rect -465 -188 -453 188
rect -419 -188 -407 188
rect -465 -200 -407 -188
rect -247 188 -189 200
rect -247 -188 -235 188
rect -201 -188 -189 188
rect -247 -200 -189 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 189 188 247 200
rect 189 -188 201 188
rect 235 -188 247 188
rect 189 -200 247 -188
rect 407 188 465 200
rect 407 -188 419 188
rect 453 -188 465 188
rect 407 -200 465 -188
<< mvndiffc >>
rect -453 -188 -419 188
rect -235 -188 -201 188
rect -17 -188 17 188
rect 201 -188 235 188
rect 419 -188 453 188
<< mvpsubdiff >>
rect -599 410 599 422
rect -599 376 -491 410
rect 491 376 599 410
rect -599 364 599 376
rect -599 314 -541 364
rect -599 -314 -587 314
rect -553 -314 -541 314
rect 541 314 599 364
rect -599 -364 -541 -314
rect 541 -314 553 314
rect 587 -314 599 314
rect 541 -364 599 -314
rect -599 -376 599 -364
rect -599 -410 -491 -376
rect 491 -410 599 -376
rect -599 -422 599 -410
<< mvpsubdiffcont >>
rect -491 376 491 410
rect -587 -314 -553 314
rect 553 -314 587 314
rect -491 -410 491 -376
<< poly >>
rect -407 272 -247 288
rect -407 238 -391 272
rect -263 238 -247 272
rect -407 200 -247 238
rect -189 272 -29 288
rect -189 238 -173 272
rect -45 238 -29 272
rect -189 200 -29 238
rect 29 272 189 288
rect 29 238 45 272
rect 173 238 189 272
rect 29 200 189 238
rect 247 272 407 288
rect 247 238 263 272
rect 391 238 407 272
rect 247 200 407 238
rect -407 -238 -247 -200
rect -407 -272 -391 -238
rect -263 -272 -247 -238
rect -407 -288 -247 -272
rect -189 -238 -29 -200
rect -189 -272 -173 -238
rect -45 -272 -29 -238
rect -189 -288 -29 -272
rect 29 -238 189 -200
rect 29 -272 45 -238
rect 173 -272 189 -238
rect 29 -288 189 -272
rect 247 -238 407 -200
rect 247 -272 263 -238
rect 391 -272 407 -238
rect 247 -288 407 -272
<< polycont >>
rect -391 238 -263 272
rect -173 238 -45 272
rect 45 238 173 272
rect 263 238 391 272
rect -391 -272 -263 -238
rect -173 -272 -45 -238
rect 45 -272 173 -238
rect 263 -272 391 -238
<< locali >>
rect -587 376 -491 410
rect 491 376 587 410
rect -587 314 -553 376
rect 553 314 587 376
rect -407 238 -391 272
rect -263 238 -247 272
rect -189 238 -173 272
rect -45 238 -29 272
rect 29 238 45 272
rect 173 238 189 272
rect 247 238 263 272
rect 391 238 407 272
rect -453 188 -419 204
rect -453 -204 -419 -188
rect -235 188 -201 204
rect -235 -204 -201 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 201 188 235 204
rect 201 -204 235 -188
rect 419 188 453 204
rect 419 -204 453 -188
rect -407 -272 -391 -238
rect -263 -272 -247 -238
rect -189 -272 -173 -238
rect -45 -272 -29 -238
rect 29 -272 45 -238
rect 173 -272 189 -238
rect 247 -272 263 -238
rect 391 -272 407 -238
rect -587 -376 -553 -314
rect 553 -376 587 -314
rect -587 -410 -491 -376
rect 491 -410 587 -376
<< viali >>
rect -391 238 -263 272
rect -173 238 -45 272
rect 45 238 173 272
rect 263 238 391 272
rect -453 -188 -419 188
rect -235 -188 -201 188
rect -17 -188 17 188
rect 201 -188 235 188
rect 419 -188 453 188
rect -391 -272 -263 -238
rect -173 -272 -45 -238
rect 45 -272 173 -238
rect 263 -272 391 -238
<< metal1 >>
rect -403 272 -251 278
rect -403 238 -391 272
rect -263 238 -251 272
rect -403 232 -251 238
rect -185 272 -33 278
rect -185 238 -173 272
rect -45 238 -33 272
rect -185 232 -33 238
rect 33 272 185 278
rect 33 238 45 272
rect 173 238 185 272
rect 33 232 185 238
rect 251 272 403 278
rect 251 238 263 272
rect 391 238 403 272
rect 251 232 403 238
rect -459 188 -413 200
rect -459 -188 -453 188
rect -419 -188 -413 188
rect -459 -200 -413 -188
rect -241 188 -195 200
rect -241 -188 -235 188
rect -201 -188 -195 188
rect -241 -200 -195 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 195 188 241 200
rect 195 -188 201 188
rect 235 -188 241 188
rect 195 -200 241 -188
rect 413 188 459 200
rect 413 -188 419 188
rect 453 -188 459 188
rect 413 -200 459 -188
rect -403 -238 -251 -232
rect -403 -272 -391 -238
rect -263 -272 -251 -238
rect -403 -278 -251 -272
rect -185 -238 -33 -232
rect -185 -272 -173 -238
rect -45 -272 -33 -238
rect -185 -278 -33 -272
rect 33 -238 185 -232
rect 33 -272 45 -238
rect 173 -272 185 -238
rect 33 -278 185 -272
rect 251 -238 403 -232
rect 251 -272 263 -238
rect 391 -272 403 -238
rect 251 -278 403 -272
<< properties >>
string FIXED_BBOX -570 -393 570 393
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2.0 l 0.8 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
