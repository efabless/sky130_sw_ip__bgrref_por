magic
tech sky130A
magscale 1 2
timestamp 1717527227
<< locali >>
rect 26884 -291054 28528 -291024
rect 26884 -291092 27004 -291054
rect 28410 -291092 28528 -291054
rect 26884 -291100 28528 -291092
rect 26884 -291994 26906 -291100
rect 26944 -291108 28528 -291100
rect 26944 -291146 28456 -291108
rect 26944 -291994 26990 -291146
rect 26884 -292046 26990 -291994
rect 28422 -292002 28456 -291146
rect 28494 -292002 28528 -291108
rect 28422 -292040 28528 -292002
rect 26892 -292244 26998 -292216
rect 26892 -292784 26924 -292244
rect 26966 -292784 26998 -292244
rect 26892 -292802 26998 -292784
rect 28422 -292274 28528 -292210
rect 28422 -292802 28460 -292274
rect 26892 -292814 28460 -292802
rect 28502 -292814 28528 -292274
rect 26892 -292860 28528 -292814
rect 26892 -292898 27040 -292860
rect 28446 -292898 28528 -292860
rect 26892 -292924 28528 -292898
<< viali >>
rect 27004 -291092 28410 -291054
rect 26906 -291994 26944 -291100
rect 28456 -292002 28494 -291108
rect 26924 -292784 26966 -292244
rect 28460 -292814 28502 -292274
rect 27040 -292898 28446 -292860
<< metal1 >>
rect 26884 -291054 28528 -291024
rect 26884 -291092 27004 -291054
rect 28410 -291092 28528 -291054
rect 26884 -291100 28528 -291092
rect 26884 -291994 26906 -291100
rect 26944 -291108 28528 -291100
rect 26944 -291146 28456 -291108
rect 26944 -291994 26990 -291146
rect 26884 -292046 26990 -291994
rect 27160 -292024 27194 -291250
rect 27320 -292024 27354 -291252
rect 27062 -292108 27354 -292024
rect 26892 -292244 26998 -292216
rect 26892 -292784 26924 -292244
rect 26966 -292784 26998 -292244
rect 27160 -292694 27194 -292108
rect 27320 -292696 27354 -292108
rect 27420 -292014 27512 -291890
rect 27748 -292014 27782 -291252
rect 27908 -292014 27942 -291252
rect 28066 -292014 28100 -291252
rect 28224 -292014 28258 -291250
rect 27420 -292096 28258 -292014
rect 28422 -292002 28456 -291146
rect 28494 -292002 28528 -291108
rect 28422 -292040 28528 -292002
rect 27420 -292186 27512 -292096
rect 27748 -292696 27782 -292096
rect 27908 -292696 27942 -292096
rect 28066 -292696 28100 -292096
rect 28224 -292694 28258 -292096
rect 28422 -292274 28528 -292210
rect 26892 -292802 26998 -292784
rect 28422 -292802 28460 -292274
rect 26892 -292814 28460 -292802
rect 28502 -292814 28528 -292274
rect 26892 -292860 28528 -292814
rect 26892 -292898 27040 -292860
rect 28446 -292898 28528 -292860
rect 26892 -292924 28528 -292898
<< metal2 >>
rect 26862 -291518 28544 -291236
rect 28470 -291608 28556 -291606
rect 26964 -291890 27512 -291608
rect 27646 -291890 28556 -291608
rect 26866 -292108 27194 -292024
rect 27420 -292186 27512 -291890
rect 28470 -292186 28556 -291890
rect 26960 -292468 27512 -292186
rect 27646 -292464 28556 -292186
rect 27646 -292468 28550 -292464
rect 26880 -292878 28562 -292616
use por_via_2cut  por_via_2cut_0
timestamp 1717527227
transform 0 1 34868 -1 0 -276416
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_1
timestamp 1717527227
transform 0 1 36220 -1 0 -276339
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_2
timestamp 1717527227
transform 0 1 35903 -1 0 -276340
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_3
timestamp 1717527227
transform 0 1 35585 -1 0 -276340
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_4
timestamp 1717527227
transform 0 1 35318 -1 0 -276340
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_5
timestamp 1717527227
transform 0 1 34996 -1 0 -276341
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_6
timestamp 1717527227
transform 0 1 35162 -1 0 -276410
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_7
timestamp 1717527227
transform 0 1 35742 -1 0 -276410
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_8
timestamp 1717527227
transform 0 1 36062 -1 0 -276408
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_9
timestamp 1717527227
transform 0 1 36356 -1 0 -276422
box 16088 -7932 16222 -7868
use por_via_4cut  por_via_4cut_0
timestamp 1717527227
transform 0 1 35160 -1 0 -275602
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_1
timestamp 1717527227
transform -1 0 43288 0 -1 -299966
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_5
timestamp 1717527227
transform 0 1 34866 -1 0 -275292
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_6
timestamp 1717527227
transform 0 1 35902 -1 0 -275362
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_7
timestamp 1717527227
transform 0 1 35580 -1 0 -275360
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_8
timestamp 1717527227
transform 0 1 35316 -1 0 -275360
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_9
timestamp 1717527227
transform 0 1 35000 -1 0 -275362
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_10
timestamp 1717527227
transform -1 0 43652 0 -1 -299954
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_14
timestamp 1717527227
transform 0 1 36058 -1 0 -275600
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_15
timestamp 1717527227
transform 0 1 35750 -1 0 -275604
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_16
timestamp 1717527227
transform 0 1 36224 -1 0 -275360
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_17
timestamp 1717527227
transform 0 1 36350 -1 0 -275290
box 15948 -7932 16222 -7868
use sky130_fd_pr__nfet_g5v0d10v5_X6E435  sky130_fd_pr__nfet_g5v0d10v5_X6E435_0
timestamp 1717527227
transform 1 0 27249 0 1 -292532
box -367 -358 367 358
use sky130_fd_pr__nfet_g5v0d10v5_Z6E439  sky130_fd_pr__nfet_g5v0d10v5_Z6E439_0
timestamp 1717527227
transform 1 0 28001 0 1 -292532
box -515 -358 515 358
use sky130_fd_pr__pfet_g5v0d10v5_CAF9E7  sky130_fd_pr__pfet_g5v0d10v5_CAF9E7_0
timestamp 1717527227
transform 1 0 27261 0 1 -291567
box -387 -547 387 547
use sky130_fd_pr__pfet_g5v0d10v5_CAPB68  sky130_fd_pr__pfet_g5v0d10v5_CAPB68_0
timestamp 1717527227
transform 1 0 28003 0 1 -291567
box -545 -547 545 547
<< end >>
