magic
tech sky130A
magscale 1 2
timestamp 1731433208
<< locali >>
rect 26884 -291054 28788 -291024
rect 26884 -291092 27004 -291054
rect 28670 -291092 28788 -291054
rect 26884 -291100 28788 -291092
rect 26884 -291994 26906 -291100
rect 26944 -291108 28788 -291100
rect 26944 -291146 28716 -291108
rect 26944 -291994 26990 -291146
rect 26884 -292046 26990 -291994
rect 28682 -292002 28716 -291146
rect 28754 -292002 28788 -291108
rect 28682 -292040 28788 -292002
rect 26892 -292244 26998 -292216
rect 26892 -292784 26924 -292244
rect 26966 -292784 26998 -292244
rect 26892 -292802 26998 -292784
rect 28682 -292274 28788 -292210
rect 28682 -292802 28720 -292274
rect 26892 -292814 28720 -292802
rect 28762 -292814 28788 -292274
rect 26892 -292860 28788 -292814
rect 26892 -292898 27040 -292860
rect 28706 -292898 28788 -292860
rect 26892 -292924 28788 -292898
<< viali >>
rect 27004 -291092 28670 -291054
rect 26906 -291994 26944 -291100
rect 28716 -292002 28754 -291108
rect 26924 -292784 26966 -292244
rect 28720 -292814 28762 -292274
rect 27040 -292898 28706 -292860
<< metal1 >>
rect 28162 -288871 28630 -288807
rect 28162 -288943 28226 -288871
rect 25940 -289007 28228 -288943
rect 28360 -289091 28457 -289004
rect 25940 -289188 28457 -289091
rect 25953 -289790 28470 -289693
rect 25940 -289937 28240 -289873
rect 28373 -289934 28470 -289790
rect 28174 -290000 28240 -289937
rect 28566 -290000 28630 -288871
rect 28174 -290064 28630 -290000
rect 28566 -290771 28630 -290064
rect 28547 -290772 28816 -290771
rect 28537 -290778 28816 -290772
rect 28537 -290866 28557 -290778
rect 28807 -290866 28816 -290778
rect 28537 -290875 28816 -290866
rect 26884 -291054 28788 -291024
rect 26884 -291092 27004 -291054
rect 28670 -291092 28788 -291054
rect 26884 -291100 28788 -291092
rect 26884 -291994 26906 -291100
rect 26944 -291108 28788 -291100
rect 26944 -291146 28716 -291108
rect 26944 -291994 26990 -291146
rect 26884 -292046 26990 -291994
rect 27160 -292024 27194 -291250
rect 27320 -292024 27354 -291252
rect 27062 -292108 27354 -292024
rect 26892 -292244 26998 -292216
rect 26892 -292784 26924 -292244
rect 26966 -292784 26998 -292244
rect 27160 -292694 27194 -292108
rect 27320 -292696 27354 -292108
rect 27420 -292014 27512 -291890
rect 27748 -292014 27782 -291252
rect 27908 -292014 27942 -291252
rect 28335 -292007 28363 -291240
rect 28495 -292006 28523 -291240
rect 28682 -292002 28716 -291146
rect 28754 -292002 28788 -291108
rect 28495 -292007 28549 -292006
rect 27420 -292096 27942 -292014
rect 28105 -292089 28549 -292007
rect 28682 -292040 28788 -292002
rect 27420 -292186 27512 -292096
rect 27748 -292696 27782 -292096
rect 27908 -292696 27942 -292096
rect 28363 -292699 28391 -292089
rect 28521 -292693 28549 -292089
rect 28682 -292274 28788 -292210
rect 26892 -292802 26998 -292784
rect 28682 -292802 28720 -292274
rect 26892 -292814 28720 -292802
rect 28762 -292814 28788 -292274
rect 26892 -292860 28788 -292814
rect 26892 -292898 27040 -292860
rect 28706 -292898 28788 -292860
rect 26892 -292924 28788 -292898
<< via1 >>
rect 28557 -290866 28807 -290778
<< metal2 >>
rect 28547 -290778 28816 -290771
rect 28547 -290866 28557 -290778
rect 28807 -290866 28816 -290778
rect 28547 -290875 28816 -290866
rect 26862 -291518 28622 -291236
rect 28730 -291608 28816 -290875
rect 26964 -291890 27512 -291608
rect 27646 -291890 28039 -291608
rect 28281 -291890 28816 -291608
rect 26866 -292108 27194 -292024
rect 27420 -292186 27512 -291890
rect 27954 -292004 28037 -291890
rect 27954 -292089 28397 -292004
rect 27954 -292186 28037 -292089
rect 28730 -292186 28816 -291890
rect 26960 -292468 27512 -292186
rect 27646 -292468 28039 -292186
rect 28270 -292464 28816 -292186
rect 28270 -292468 28810 -292464
rect 26880 -292878 28822 -292616
use por_via_2cut  por_via_2cut_0
timestamp 1718283729
transform 0 1 34868 -1 0 -276416
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_1
timestamp 1718283729
transform 0 1 36200 -1 0 -276341
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_2
timestamp 1718283729
transform 0 1 35903 -1 0 -276340
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_3
timestamp 1718283729
transform 0 1 35585 -1 0 -276340
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_4
timestamp 1718283729
transform 0 1 35318 -1 0 -276340
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_5
timestamp 1718283729
transform 0 1 34996 -1 0 -276341
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_6
timestamp 1718283729
transform 0 1 35162 -1 0 -276410
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_7
timestamp 1718283729
transform 0 1 35742 -1 0 -276410
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_8
timestamp 1718283729
transform 0 1 36514 -1 0 -276343
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_9
timestamp 1718283729
transform 0 1 36354 -1 0 -276412
box 16088 -7932 16222 -7868
use por_via_4cut  por_via_4cut_0
timestamp 1718283729
transform 0 1 35160 -1 0 -275602
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_1
timestamp 1718283729
transform -1 0 43288 0 -1 -299966
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_2
timestamp 1718283729
transform 0 1 36173 -1 0 -275358
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_3
timestamp 1718283729
transform 0 1 36488 -1 0 -275363
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_4
timestamp 1718283729
transform -1 0 44336 0 -1 -299946
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_5
timestamp 1718283729
transform 0 1 34866 -1 0 -275292
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_6
timestamp 1718283729
transform 0 1 35902 -1 0 -275362
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_7
timestamp 1718283729
transform 0 1 35580 -1 0 -275360
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_8
timestamp 1718283729
transform 0 1 35316 -1 0 -275360
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_9
timestamp 1718283729
transform 0 1 35000 -1 0 -275362
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_10
timestamp 1718283729
transform -1 0 43652 0 -1 -299954
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_15
timestamp 1718283729
transform 0 1 35750 -1 0 -275604
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_16
timestamp 1718283729
transform 0 1 36325 -1 0 -275594
box 15948 -7932 16222 -7868
use sky130_fd_pr__nfet_g5v0d10v5_X6E435  sky130_fd_pr__nfet_g5v0d10v5_X6E435_0 paramcells
timestamp 1718283729
transform 1 0 27249 0 1 -292532
box -367 -358 367 358
use sky130_fd_pr__nfet_g5v0d10v5_X6E435  sky130_fd_pr__nfet_g5v0d10v5_X6E435_1
timestamp 1718283729
transform 1 0 27853 0 1 -292532
box -367 -358 367 358
use sky130_fd_pr__nfet_g5v0d10v5_X6E435  sky130_fd_pr__nfet_g5v0d10v5_X6E435_2
timestamp 1718283729
transform 1 0 28457 0 1 -292532
box -367 -358 367 358
use sky130_fd_pr__pfet_g5v0d10v5_CAF9E7  sky130_fd_pr__pfet_g5v0d10v5_CAF9E7_0 paramcells
timestamp 1718283729
transform 1 0 27845 0 1 -291567
box -387 -547 387 547
use sky130_fd_pr__pfet_g5v0d10v5_CAF9E7  sky130_fd_pr__pfet_g5v0d10v5_CAF9E7_1
timestamp 1718283729
transform 1 0 27261 0 1 -291567
box -387 -547 387 547
use sky130_fd_pr__pfet_g5v0d10v5_CAF9E7  sky130_fd_pr__pfet_g5v0d10v5_CAF9E7_2
timestamp 1718283729
transform 1 0 28429 0 1 -291567
box -387 -547 387 547
use sky130_fd_sc_hvl__inv_16  sky130_fd_sc_hvl__inv_16_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1729530005
transform 1 0 25658 0 -1 -288632
box -66 -43 2754 897
use sky130_fd_sc_hvl__inv_16  sky130_fd_sc_hvl__inv_16_1
timestamp 1729530005
transform 1 0 25658 0 1 -290260
box -66 -43 2754 897
<< end >>
