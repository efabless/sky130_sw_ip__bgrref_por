magic
tech sky130A
magscale 1 2
timestamp 1717527227
<< nwell >>
rect -545 -547 545 547
<< mvpmos >>
rect -287 -250 -187 250
rect -129 -250 -29 250
rect 29 -250 129 250
rect 187 -250 287 250
<< mvpdiff >>
rect -345 238 -287 250
rect -345 -238 -333 238
rect -299 -238 -287 238
rect -345 -250 -287 -238
rect -187 238 -129 250
rect -187 -238 -175 238
rect -141 -238 -129 238
rect -187 -250 -129 -238
rect -29 238 29 250
rect -29 -238 -17 238
rect 17 -238 29 238
rect -29 -250 29 -238
rect 129 238 187 250
rect 129 -238 141 238
rect 175 -238 187 238
rect 129 -250 187 -238
rect 287 238 345 250
rect 287 -238 299 238
rect 333 -238 345 238
rect 287 -250 345 -238
<< mvpdiffc >>
rect -333 -238 -299 238
rect -175 -238 -141 238
rect -17 -238 17 238
rect 141 -238 175 238
rect 299 -238 333 238
<< mvnsubdiff >>
rect -479 469 479 481
rect -479 435 -371 469
rect 371 435 479 469
rect -479 423 479 435
rect -479 373 -421 423
rect -479 -373 -467 373
rect -433 -373 -421 373
rect 421 373 479 423
rect -479 -423 -421 -373
rect 421 -373 433 373
rect 467 -373 479 373
rect 421 -423 479 -373
rect -479 -435 479 -423
rect -479 -469 -371 -435
rect 371 -469 479 -435
rect -479 -481 479 -469
<< mvnsubdiffcont >>
rect -371 435 371 469
rect -467 -373 -433 373
rect 433 -373 467 373
rect -371 -469 371 -435
<< poly >>
rect -287 331 -187 347
rect -287 297 -271 331
rect -203 297 -187 331
rect -287 250 -187 297
rect -129 331 -29 347
rect -129 297 -113 331
rect -45 297 -29 331
rect -129 250 -29 297
rect 29 331 129 347
rect 29 297 45 331
rect 113 297 129 331
rect 29 250 129 297
rect 187 331 287 347
rect 187 297 203 331
rect 271 297 287 331
rect 187 250 287 297
rect -287 -297 -187 -250
rect -287 -331 -271 -297
rect -203 -331 -187 -297
rect -287 -347 -187 -331
rect -129 -297 -29 -250
rect -129 -331 -113 -297
rect -45 -331 -29 -297
rect -129 -347 -29 -331
rect 29 -297 129 -250
rect 29 -331 45 -297
rect 113 -331 129 -297
rect 29 -347 129 -331
rect 187 -297 287 -250
rect 187 -331 203 -297
rect 271 -331 287 -297
rect 187 -347 287 -331
<< polycont >>
rect -271 297 -203 331
rect -113 297 -45 331
rect 45 297 113 331
rect 203 297 271 331
rect -271 -331 -203 -297
rect -113 -331 -45 -297
rect 45 -331 113 -297
rect 203 -331 271 -297
<< locali >>
rect -467 435 -371 469
rect 371 435 467 469
rect -467 373 -433 435
rect 433 373 467 435
rect -287 297 -271 331
rect -203 297 -187 331
rect -129 297 -113 331
rect -45 297 -29 331
rect 29 297 45 331
rect 113 297 129 331
rect 187 297 203 331
rect 271 297 287 331
rect -333 238 -299 254
rect -333 -254 -299 -238
rect -175 238 -141 254
rect -175 -254 -141 -238
rect -17 238 17 254
rect -17 -254 17 -238
rect 141 238 175 254
rect 141 -254 175 -238
rect 299 238 333 254
rect 299 -254 333 -238
rect -287 -331 -271 -297
rect -203 -331 -187 -297
rect -129 -331 -113 -297
rect -45 -331 -29 -297
rect 29 -331 45 -297
rect 113 -331 129 -297
rect 187 -331 203 -297
rect 271 -331 287 -297
rect -467 -435 -433 -373
rect 433 -435 467 -373
rect -467 -469 -371 -435
rect 371 -469 467 -435
<< viali >>
rect -271 297 -203 331
rect -113 297 -45 331
rect 45 297 113 331
rect 203 297 271 331
rect -333 -238 -299 238
rect -175 -238 -141 238
rect -17 -238 17 238
rect 141 -238 175 238
rect 299 -238 333 238
rect -271 -331 -203 -297
rect -113 -331 -45 -297
rect 45 -331 113 -297
rect 203 -331 271 -297
<< metal1 >>
rect -283 331 -191 337
rect -283 297 -271 331
rect -203 297 -191 331
rect -283 291 -191 297
rect -125 331 -33 337
rect -125 297 -113 331
rect -45 297 -33 331
rect -125 291 -33 297
rect 33 331 125 337
rect 33 297 45 331
rect 113 297 125 331
rect 33 291 125 297
rect 191 331 283 337
rect 191 297 203 331
rect 271 297 283 331
rect 191 291 283 297
rect -339 238 -293 250
rect -339 -238 -333 238
rect -299 -238 -293 238
rect -339 -250 -293 -238
rect -181 238 -135 250
rect -181 -238 -175 238
rect -141 -238 -135 238
rect -181 -250 -135 -238
rect -23 238 23 250
rect -23 -238 -17 238
rect 17 -238 23 238
rect -23 -250 23 -238
rect 135 238 181 250
rect 135 -238 141 238
rect 175 -238 181 238
rect 135 -250 181 -238
rect 293 238 339 250
rect 293 -238 299 238
rect 333 -238 339 238
rect 293 -250 339 -238
rect -283 -297 -191 -291
rect -283 -331 -271 -297
rect -203 -331 -191 -297
rect -283 -337 -191 -331
rect -125 -297 -33 -291
rect -125 -331 -113 -297
rect -45 -331 -33 -297
rect -125 -337 -33 -331
rect 33 -297 125 -291
rect 33 -331 45 -297
rect 113 -331 125 -297
rect 33 -337 125 -331
rect 191 -297 283 -291
rect 191 -331 203 -297
rect 271 -331 283 -297
rect 191 -337 283 -331
<< properties >>
string FIXED_BBOX -450 -452 450 452
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2.5 l 0.50 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
