magic
tech sky130A
magscale 1 2
timestamp 1717527330
<< metal3 >>
rect -17940 3472 -14468 3500
rect -17940 448 -14552 3472
rect -14488 448 -14468 3472
rect -17940 420 -14468 448
rect -13642 3472 -10170 3500
rect -13642 448 -10254 3472
rect -10190 448 -10170 3472
rect -13642 420 -10170 448
rect -9344 3472 -5872 3500
rect -9344 448 -5956 3472
rect -5892 448 -5872 3472
rect -9344 420 -5872 448
rect -5046 3472 -1574 3500
rect -5046 448 -1658 3472
rect -1594 448 -1574 3472
rect -5046 420 -1574 448
rect -748 3472 2724 3500
rect -748 448 2640 3472
rect 2704 448 2724 3472
rect -748 420 2724 448
rect 3550 3472 7022 3500
rect 3550 448 6938 3472
rect 7002 448 7022 3472
rect 3550 420 7022 448
rect 7848 3472 11320 3500
rect 7848 448 11236 3472
rect 11300 448 11320 3472
rect 7848 420 11320 448
rect 12146 3472 15618 3500
rect 12146 448 15534 3472
rect 15598 448 15618 3472
rect 12146 420 15618 448
rect 16444 3472 19916 3500
rect 16444 448 19832 3472
rect 19896 448 19916 3472
rect 16444 420 19916 448
rect 20742 3472 24214 3500
rect 20742 448 24130 3472
rect 24194 448 24214 3472
rect 20742 420 24214 448
rect -17940 -148 -14468 -120
rect -17940 -3172 -14552 -148
rect -14488 -3172 -14468 -148
rect -17940 -3200 -14468 -3172
rect -13642 -148 -10170 -120
rect -13642 -3172 -10254 -148
rect -10190 -3172 -10170 -148
rect -13642 -3200 -10170 -3172
rect -9344 -148 -5872 -120
rect -9344 -3172 -5956 -148
rect -5892 -3172 -5872 -148
rect -9344 -3200 -5872 -3172
rect -5046 -148 -1574 -120
rect -5046 -3172 -1658 -148
rect -1594 -3172 -1574 -148
rect -5046 -3200 -1574 -3172
rect -748 -148 2724 -120
rect -748 -3172 2640 -148
rect 2704 -3172 2724 -148
rect -748 -3200 2724 -3172
rect 3550 -148 7022 -120
rect 3550 -3172 6938 -148
rect 7002 -3172 7022 -148
rect 3550 -3200 7022 -3172
rect 7848 -148 11320 -120
rect 7848 -3172 11236 -148
rect 11300 -3172 11320 -148
rect 7848 -3200 11320 -3172
rect 12146 -148 15618 -120
rect 12146 -3172 15534 -148
rect 15598 -3172 15618 -148
rect 12146 -3200 15618 -3172
rect 16444 -148 19916 -120
rect 16444 -3172 19832 -148
rect 19896 -3172 19916 -148
rect 16444 -3200 19916 -3172
rect 20742 -148 24214 -120
rect 20742 -3172 24130 -148
rect 24194 -3172 24214 -148
rect 20742 -3200 24214 -3172
<< via3 >>
rect -14552 448 -14488 3472
rect -10254 448 -10190 3472
rect -5956 448 -5892 3472
rect -1658 448 -1594 3472
rect 2640 448 2704 3472
rect 6938 448 7002 3472
rect 11236 448 11300 3472
rect 15534 448 15598 3472
rect 19832 448 19896 3472
rect 24130 448 24194 3472
rect -14552 -3172 -14488 -148
rect -10254 -3172 -10190 -148
rect -5956 -3172 -5892 -148
rect -1658 -3172 -1594 -148
rect 2640 -3172 2704 -148
rect 6938 -3172 7002 -148
rect 11236 -3172 11300 -148
rect 15534 -3172 15598 -148
rect 19832 -3172 19896 -148
rect 24130 -3172 24194 -148
<< mimcap >>
rect -17900 3420 -14900 3460
rect -17900 500 -17860 3420
rect -14940 500 -14900 3420
rect -17900 460 -14900 500
rect -13602 3420 -10602 3460
rect -13602 500 -13562 3420
rect -10642 500 -10602 3420
rect -13602 460 -10602 500
rect -9304 3420 -6304 3460
rect -9304 500 -9264 3420
rect -6344 500 -6304 3420
rect -9304 460 -6304 500
rect -5006 3420 -2006 3460
rect -5006 500 -4966 3420
rect -2046 500 -2006 3420
rect -5006 460 -2006 500
rect -708 3420 2292 3460
rect -708 500 -668 3420
rect 2252 500 2292 3420
rect -708 460 2292 500
rect 3590 3420 6590 3460
rect 3590 500 3630 3420
rect 6550 500 6590 3420
rect 3590 460 6590 500
rect 7888 3420 10888 3460
rect 7888 500 7928 3420
rect 10848 500 10888 3420
rect 7888 460 10888 500
rect 12186 3420 15186 3460
rect 12186 500 12226 3420
rect 15146 500 15186 3420
rect 12186 460 15186 500
rect 16484 3420 19484 3460
rect 16484 500 16524 3420
rect 19444 500 19484 3420
rect 16484 460 19484 500
rect 20782 3420 23782 3460
rect 20782 500 20822 3420
rect 23742 500 23782 3420
rect 20782 460 23782 500
rect -17900 -200 -14900 -160
rect -17900 -3120 -17860 -200
rect -14940 -3120 -14900 -200
rect -17900 -3160 -14900 -3120
rect -13602 -200 -10602 -160
rect -13602 -3120 -13562 -200
rect -10642 -3120 -10602 -200
rect -13602 -3160 -10602 -3120
rect -9304 -200 -6304 -160
rect -9304 -3120 -9264 -200
rect -6344 -3120 -6304 -200
rect -9304 -3160 -6304 -3120
rect -5006 -200 -2006 -160
rect -5006 -3120 -4966 -200
rect -2046 -3120 -2006 -200
rect -5006 -3160 -2006 -3120
rect -708 -200 2292 -160
rect -708 -3120 -668 -200
rect 2252 -3120 2292 -200
rect -708 -3160 2292 -3120
rect 3590 -200 6590 -160
rect 3590 -3120 3630 -200
rect 6550 -3120 6590 -200
rect 3590 -3160 6590 -3120
rect 7888 -200 10888 -160
rect 7888 -3120 7928 -200
rect 10848 -3120 10888 -200
rect 7888 -3160 10888 -3120
rect 12186 -200 15186 -160
rect 12186 -3120 12226 -200
rect 15146 -3120 15186 -200
rect 12186 -3160 15186 -3120
rect 16484 -200 19484 -160
rect 16484 -3120 16524 -200
rect 19444 -3120 19484 -200
rect 16484 -3160 19484 -3120
rect 20782 -200 23782 -160
rect 20782 -3120 20822 -200
rect 23742 -3120 23782 -200
rect 20782 -3160 23782 -3120
<< mimcapcontact >>
rect -17860 500 -14940 3420
rect -13562 500 -10642 3420
rect -9264 500 -6344 3420
rect -4966 500 -2046 3420
rect -668 500 2252 3420
rect 3630 500 6550 3420
rect 7928 500 10848 3420
rect 12226 500 15146 3420
rect 16524 500 19444 3420
rect 20822 500 23742 3420
rect -17860 -3120 -14940 -200
rect -13562 -3120 -10642 -200
rect -9264 -3120 -6344 -200
rect -4966 -3120 -2046 -200
rect -668 -3120 2252 -200
rect 3630 -3120 6550 -200
rect 7928 -3120 10848 -200
rect 12226 -3120 15146 -200
rect 16524 -3120 19444 -200
rect 20822 -3120 23742 -200
<< metal4 >>
rect -16452 3421 -16348 3620
rect -14572 3472 -14468 3620
rect -17861 3420 -14939 3421
rect -17861 500 -17860 3420
rect -14940 500 -14939 3420
rect -17861 499 -14939 500
rect -16452 -199 -16348 499
rect -14572 448 -14552 3472
rect -14488 448 -14468 3472
rect -12154 3421 -12050 3620
rect -10274 3472 -10170 3620
rect -13563 3420 -10641 3421
rect -13563 500 -13562 3420
rect -10642 500 -10641 3420
rect -13563 499 -10641 500
rect -14572 -148 -14468 448
rect -17861 -200 -14939 -199
rect -17861 -3120 -17860 -200
rect -14940 -3120 -14939 -200
rect -17861 -3121 -14939 -3120
rect -16452 -3320 -16348 -3121
rect -14572 -3172 -14552 -148
rect -14488 -3172 -14468 -148
rect -12154 -199 -12050 499
rect -10274 448 -10254 3472
rect -10190 448 -10170 3472
rect -7856 3421 -7752 3620
rect -5976 3472 -5872 3620
rect -9265 3420 -6343 3421
rect -9265 500 -9264 3420
rect -6344 500 -6343 3420
rect -9265 499 -6343 500
rect -10274 -148 -10170 448
rect -13563 -200 -10641 -199
rect -13563 -3120 -13562 -200
rect -10642 -3120 -10641 -200
rect -13563 -3121 -10641 -3120
rect -14572 -3320 -14468 -3172
rect -12154 -3320 -12050 -3121
rect -10274 -3172 -10254 -148
rect -10190 -3172 -10170 -148
rect -7856 -199 -7752 499
rect -5976 448 -5956 3472
rect -5892 448 -5872 3472
rect -3558 3421 -3454 3620
rect -1678 3472 -1574 3620
rect -4967 3420 -2045 3421
rect -4967 500 -4966 3420
rect -2046 500 -2045 3420
rect -4967 499 -2045 500
rect -5976 -148 -5872 448
rect -9265 -200 -6343 -199
rect -9265 -3120 -9264 -200
rect -6344 -3120 -6343 -200
rect -9265 -3121 -6343 -3120
rect -10274 -3320 -10170 -3172
rect -7856 -3320 -7752 -3121
rect -5976 -3172 -5956 -148
rect -5892 -3172 -5872 -148
rect -3558 -199 -3454 499
rect -1678 448 -1658 3472
rect -1594 448 -1574 3472
rect 740 3421 844 3620
rect 2620 3472 2724 3620
rect -669 3420 2253 3421
rect -669 500 -668 3420
rect 2252 500 2253 3420
rect -669 499 2253 500
rect -1678 -148 -1574 448
rect -4967 -200 -2045 -199
rect -4967 -3120 -4966 -200
rect -2046 -3120 -2045 -200
rect -4967 -3121 -2045 -3120
rect -5976 -3320 -5872 -3172
rect -3558 -3320 -3454 -3121
rect -1678 -3172 -1658 -148
rect -1594 -3172 -1574 -148
rect 740 -199 844 499
rect 2620 448 2640 3472
rect 2704 448 2724 3472
rect 5038 3421 5142 3620
rect 6918 3472 7022 3620
rect 3629 3420 6551 3421
rect 3629 500 3630 3420
rect 6550 500 6551 3420
rect 3629 499 6551 500
rect 2620 -148 2724 448
rect -669 -200 2253 -199
rect -669 -3120 -668 -200
rect 2252 -3120 2253 -200
rect -669 -3121 2253 -3120
rect -1678 -3320 -1574 -3172
rect 740 -3320 844 -3121
rect 2620 -3172 2640 -148
rect 2704 -3172 2724 -148
rect 5038 -199 5142 499
rect 6918 448 6938 3472
rect 7002 448 7022 3472
rect 9336 3421 9440 3620
rect 11216 3472 11320 3620
rect 7927 3420 10849 3421
rect 7927 500 7928 3420
rect 10848 500 10849 3420
rect 7927 499 10849 500
rect 6918 -148 7022 448
rect 3629 -200 6551 -199
rect 3629 -3120 3630 -200
rect 6550 -3120 6551 -200
rect 3629 -3121 6551 -3120
rect 2620 -3320 2724 -3172
rect 5038 -3320 5142 -3121
rect 6918 -3172 6938 -148
rect 7002 -3172 7022 -148
rect 9336 -199 9440 499
rect 11216 448 11236 3472
rect 11300 448 11320 3472
rect 13634 3421 13738 3620
rect 15514 3472 15618 3620
rect 12225 3420 15147 3421
rect 12225 500 12226 3420
rect 15146 500 15147 3420
rect 12225 499 15147 500
rect 11216 -148 11320 448
rect 7927 -200 10849 -199
rect 7927 -3120 7928 -200
rect 10848 -3120 10849 -200
rect 7927 -3121 10849 -3120
rect 6918 -3320 7022 -3172
rect 9336 -3320 9440 -3121
rect 11216 -3172 11236 -148
rect 11300 -3172 11320 -148
rect 13634 -199 13738 499
rect 15514 448 15534 3472
rect 15598 448 15618 3472
rect 17932 3421 18036 3620
rect 19812 3472 19916 3620
rect 16523 3420 19445 3421
rect 16523 500 16524 3420
rect 19444 500 19445 3420
rect 16523 499 19445 500
rect 15514 -148 15618 448
rect 12225 -200 15147 -199
rect 12225 -3120 12226 -200
rect 15146 -3120 15147 -200
rect 12225 -3121 15147 -3120
rect 11216 -3320 11320 -3172
rect 13634 -3320 13738 -3121
rect 15514 -3172 15534 -148
rect 15598 -3172 15618 -148
rect 17932 -199 18036 499
rect 19812 448 19832 3472
rect 19896 448 19916 3472
rect 22230 3421 22334 3620
rect 24110 3472 24214 3620
rect 20821 3420 23743 3421
rect 20821 500 20822 3420
rect 23742 500 23743 3420
rect 20821 499 23743 500
rect 19812 -148 19916 448
rect 16523 -200 19445 -199
rect 16523 -3120 16524 -200
rect 19444 -3120 19445 -200
rect 16523 -3121 19445 -3120
rect 15514 -3320 15618 -3172
rect 17932 -3320 18036 -3121
rect 19812 -3172 19832 -148
rect 19896 -3172 19916 -148
rect 22230 -199 22334 499
rect 24110 448 24130 3472
rect 24194 448 24214 3472
rect 24110 -148 24214 448
rect 20821 -200 23743 -199
rect 20821 -3120 20822 -200
rect 23742 -3120 23743 -200
rect 20821 -3121 23743 -3120
rect 19812 -3320 19916 -3172
rect 22230 -3320 22334 -3121
rect 24110 -3172 24130 -148
rect 24194 -3172 24214 -148
rect 24110 -3320 24214 -3172
<< properties >>
string FIXED_BBOX 14568 120 17648 3200
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 15.00 l 15.00 val 461.4 carea 2.00 cperi 0.19 nx 10 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
