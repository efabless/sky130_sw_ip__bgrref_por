magic
tech sky130A
magscale 1 2
timestamp 1717613630
<< pwell >>
rect 28622 -284511 28714 -284488
<< locali >>
rect 22374 -282879 22595 -282768
rect 22374 -285902 22449 -282879
rect 16607 -285909 22449 -285902
rect 22500 -285909 22595 -282879
rect 23106 -283911 25430 -283880
rect 23106 -283964 23154 -283911
rect 25400 -283964 25430 -283911
rect 23106 -284014 25430 -283964
rect 28622 -284463 28714 -284449
rect 28622 -284507 28637 -284463
rect 28698 -284507 28714 -284463
rect 28622 -284521 28714 -284507
rect 23927 -285574 25419 -285456
rect 23927 -285576 23981 -285574
rect 23224 -285638 23981 -285576
rect 24303 -285638 24413 -285574
rect 25378 -285638 25419 -285574
rect 23224 -285668 25419 -285638
rect 23927 -285670 25419 -285668
rect 16607 -285970 22595 -285909
rect 16607 -286004 22591 -285970
rect 16617 -286412 22601 -286310
rect 26242 -286341 30542 -286311
rect 22968 -286380 25227 -286367
rect 22968 -286430 23073 -286380
rect 25187 -286430 25227 -286380
rect 26242 -286392 26290 -286341
rect 30511 -286392 30542 -286341
rect 26242 -286419 30542 -286392
rect 22968 -286523 25227 -286430
rect 31688 -286470 32882 -286441
rect 30834 -286500 31401 -286477
rect 30834 -286538 30990 -286500
rect 31307 -286531 31401 -286500
rect 31307 -286538 31346 -286531
rect 30834 -286555 31346 -286538
rect 25699 -286846 26258 -286845
rect 25699 -286880 26260 -286846
rect 25699 -286926 25738 -286880
rect 26202 -286926 26260 -286880
rect 25699 -286941 26260 -286926
rect 25705 -286943 26260 -286941
rect 22361 -287116 22514 -287045
rect 22361 -289459 22409 -287116
rect 22456 -289459 22514 -287116
rect 31325 -287471 31346 -286555
rect 31380 -287471 31401 -286531
rect 31688 -286595 31722 -286470
rect 32843 -286595 32882 -286470
rect 31688 -286651 32882 -286595
rect 31325 -287505 31401 -287471
rect 31224 -288061 32867 -288047
rect 31224 -288116 32066 -288061
rect 32836 -288116 32867 -288061
rect 31224 -288219 32867 -288116
rect 26938 -288593 30425 -288542
rect 26938 -288658 27023 -288593
rect 30391 -288658 30425 -288593
rect 26938 -288686 30425 -288658
rect 31214 -288637 32867 -288616
rect 31214 -288681 31243 -288637
rect 32843 -288681 32867 -288637
rect 31214 -288693 32867 -288681
rect 22361 -289507 22514 -289459
<< viali >>
rect 22449 -285909 22500 -282879
rect 23154 -283964 25400 -283911
rect 28637 -284507 28698 -284463
rect 27863 -284571 27973 -284536
rect 27781 -284649 27889 -284615
rect 28265 -284757 28299 -284640
rect 28374 -284645 28408 -284528
rect 30110 -284776 30161 -284624
rect 27316 -285199 27424 -285165
rect 28103 -285234 28137 -285117
rect 28370 -285212 28404 -285095
rect 30110 -285111 30161 -284959
rect 28637 -285276 28698 -285232
rect 23981 -285638 24303 -285574
rect 24413 -285638 25378 -285574
rect 23073 -286430 25187 -286380
rect 26290 -286392 30511 -286341
rect 30990 -286538 31307 -286500
rect 25738 -286926 26202 -286880
rect 22409 -289459 22456 -287116
rect 31346 -287471 31380 -286531
rect 31722 -286595 32843 -286470
rect 32066 -288116 32836 -288061
rect 27023 -288658 30391 -288593
rect 31243 -288681 32843 -288637
<< metal1 >>
rect 29108 -282710 29430 -282696
rect 22374 -282879 22595 -282768
rect 29108 -282842 29132 -282710
rect 29402 -282842 29430 -282710
rect 29108 -282864 29430 -282842
rect 16742 -283415 17114 -282983
rect 17210 -283415 17582 -282983
rect 17678 -283415 18050 -282983
rect 18146 -283415 18518 -282983
rect 18614 -283415 18986 -282983
rect 19082 -283415 19454 -282983
rect 19550 -283415 19922 -282983
rect 20018 -283415 20390 -282983
rect 20486 -283415 20858 -282983
rect 20954 -283415 21326 -282983
rect 21422 -283415 21794 -282983
rect 21890 -283415 22262 -282983
rect 22374 -283561 22449 -282879
rect 22500 -283561 22595 -282879
rect 22374 -284846 22444 -283561
rect 22515 -284846 22595 -283561
rect 22374 -285345 22449 -284846
rect 22500 -285345 22595 -284846
rect 16739 -286950 16883 -285381
rect 22374 -285383 22444 -285345
rect 16975 -285816 17349 -285384
rect 17443 -285816 17817 -285384
rect 17911 -285816 18285 -285384
rect 18379 -285816 18753 -285384
rect 18847 -285816 19221 -285384
rect 19315 -285816 19689 -285384
rect 19783 -285816 20157 -285384
rect 20251 -285816 20625 -285384
rect 20719 -285816 21093 -285384
rect 21187 -285816 21561 -285384
rect 21655 -285816 22029 -285384
rect 22124 -285816 22444 -285383
rect 22374 -285914 22444 -285816
rect 22515 -285914 22595 -285345
rect 22374 -285970 22595 -285914
rect 22729 -283158 22966 -283152
rect 22729 -285435 22966 -283451
rect 29212 -283744 29314 -282864
rect 23069 -283911 25750 -283855
rect 23069 -283964 23154 -283911
rect 25400 -283964 25750 -283911
rect 23069 -284018 25750 -283964
rect 23099 -284113 23437 -284073
rect 23568 -284112 23906 -284080
rect 24012 -284109 24232 -284076
rect 24345 -284109 24536 -284076
rect 23099 -284317 23155 -284113
rect 23099 -284357 23447 -284317
rect 23568 -284323 23600 -284112
rect 23568 -284355 23904 -284323
rect 24012 -284325 24045 -284109
rect 24345 -284325 24378 -284109
rect 24661 -284111 24868 -284078
rect 24975 -284111 25263 -284078
rect 25587 -284082 25750 -284018
rect 29212 -284040 29230 -283744
rect 29302 -284040 29314 -283744
rect 29212 -284062 29314 -284040
rect 24661 -284320 24694 -284111
rect 24975 -284316 25008 -284111
rect 25587 -284182 27265 -284082
rect 25587 -284245 30386 -284182
rect 23099 -284613 23155 -284357
rect 23018 -284682 23155 -284613
rect 22729 -286051 22740 -285435
rect 22952 -286051 22966 -285435
rect 22729 -286068 22966 -286051
rect 23099 -284697 23155 -284682
rect 23099 -284737 23434 -284697
rect 23568 -284714 23600 -284355
rect 24012 -284358 24229 -284325
rect 24345 -284358 24543 -284325
rect 24661 -284353 24866 -284320
rect 24975 -284349 25275 -284316
rect 24012 -284714 24045 -284358
rect 23099 -285026 23155 -284737
rect 23568 -284746 23781 -284714
rect 23473 -284835 23515 -284829
rect 23568 -284835 23600 -284746
rect 23473 -284957 23600 -284835
rect 23099 -285066 23431 -285026
rect 23099 -285133 23155 -285066
rect 23099 -285173 23437 -285133
rect 23099 -285479 23155 -285173
rect 23099 -285519 23444 -285479
rect 23099 -286128 23155 -285519
rect 23473 -285990 23515 -284957
rect 23568 -285044 23600 -284957
rect 24012 -284747 24212 -284714
rect 24345 -284716 24378 -284358
rect 24661 -284712 24694 -284353
rect 24012 -284985 24045 -284747
rect 24345 -284749 24549 -284716
rect 24661 -284745 24833 -284712
rect 24975 -284714 25008 -284349
rect 25619 -284540 25768 -284501
rect 24345 -284983 24378 -284749
rect 24661 -284979 24694 -284745
rect 24975 -284747 25263 -284714
rect 24975 -284974 25008 -284747
rect 24012 -285018 24222 -284985
rect 24345 -285016 24534 -284983
rect 24661 -285012 24843 -284979
rect 24975 -285007 25262 -284974
rect 23568 -285076 23775 -285044
rect 23568 -285153 23600 -285076
rect 24012 -285089 24045 -285018
rect 24345 -285087 24378 -285016
rect 24661 -285087 24694 -285012
rect 24012 -285122 24215 -285089
rect 24345 -285120 24515 -285087
rect 24661 -285120 24843 -285087
rect 24975 -285092 25008 -285007
rect 23568 -285185 23794 -285153
rect 23568 -285469 23600 -285185
rect 23568 -285501 23783 -285469
rect 23568 -285504 23600 -285501
rect 23819 -285909 23858 -285232
rect 24012 -285356 24045 -285122
rect 24012 -285389 24205 -285356
rect 24345 -285358 24378 -285120
rect 24345 -285391 24517 -285358
rect 24661 -285359 24694 -285120
rect 24975 -285125 25260 -285092
rect 24975 -285352 25008 -285125
rect 23927 -285574 24311 -285456
rect 23927 -285638 23981 -285574
rect 24303 -285638 24311 -285574
rect 23927 -285670 24311 -285638
rect 24345 -285788 24378 -285391
rect 24661 -285392 24849 -285359
rect 24975 -285385 25270 -285352
rect 24975 -285391 25008 -285385
rect 24661 -285409 24694 -285392
rect 24406 -285574 25419 -285456
rect 24406 -285638 24413 -285574
rect 25378 -285638 25419 -285574
rect 24406 -285670 25419 -285638
rect 25729 -285727 25768 -284540
rect 26002 -285371 26165 -284245
rect 26848 -284822 26944 -284333
rect 27088 -284345 30386 -284245
rect 27097 -284449 28713 -284442
rect 27097 -284463 28714 -284449
rect 27097 -284474 28637 -284463
rect 28622 -284507 28637 -284474
rect 28698 -284507 28714 -284463
rect 28367 -284528 28416 -284514
rect 28622 -284521 28714 -284507
rect 31301 -284480 31437 -284440
rect 27849 -284536 27989 -284528
rect 27849 -284571 27863 -284536
rect 27973 -284571 27989 -284536
rect 27849 -284580 27989 -284571
rect 27769 -284615 27901 -284608
rect 27769 -284649 27781 -284615
rect 27889 -284649 27901 -284615
rect 27769 -284656 27901 -284649
rect 28258 -284640 28307 -284622
rect 28258 -284757 28265 -284640
rect 28299 -284757 28307 -284640
rect 28367 -284645 28374 -284528
rect 28408 -284645 28416 -284528
rect 28367 -284662 28416 -284645
rect 30098 -284624 30174 -284613
rect 28258 -284777 28307 -284757
rect 30098 -284776 30110 -284624
rect 30161 -284670 30174 -284624
rect 31301 -284670 31341 -284480
rect 30161 -284710 31341 -284670
rect 30161 -284776 30174 -284710
rect 30098 -284790 30174 -284776
rect 26848 -284918 27244 -284822
rect 30259 -284917 30440 -284822
rect 30742 -284917 30748 -284822
rect 30098 -284959 30174 -284948
rect 28362 -285095 28412 -285078
rect 28094 -285117 28144 -285102
rect 27301 -285165 27442 -285155
rect 27301 -285199 27316 -285165
rect 27424 -285199 27442 -285165
rect 27301 -285207 27442 -285199
rect 28094 -285234 28103 -285117
rect 28137 -285234 28144 -285117
rect 28145 -285185 28151 -285150
rect 28280 -285185 28286 -285150
rect 28362 -285212 28370 -285095
rect 28404 -285212 28412 -285095
rect 30098 -285111 30110 -284959
rect 30161 -285003 30174 -284959
rect 30161 -285043 31241 -285003
rect 30161 -285111 30174 -285043
rect 30098 -285125 30174 -285111
rect 28362 -285230 28412 -285212
rect 30846 -285182 31152 -285171
rect 28094 -285254 28144 -285234
rect 28622 -285232 28714 -285218
rect 28622 -285276 28637 -285232
rect 28698 -285276 28714 -285232
rect 28622 -285291 28714 -285276
rect 30846 -285371 30857 -285182
rect 26002 -285527 30857 -285371
rect 31138 -285527 31152 -285182
rect 26002 -285534 31152 -285527
rect 27543 -285616 30899 -285577
rect 27543 -285687 30799 -285652
rect 25729 -285766 30012 -285727
rect 23929 -285798 24465 -285788
rect 23929 -285855 23949 -285798
rect 24451 -285855 24465 -285798
rect 23929 -285869 24465 -285855
rect 25576 -285848 30012 -285809
rect 25576 -285909 25615 -285848
rect 23819 -285948 25615 -285909
rect 29447 -285927 30698 -285913
rect 29225 -285960 30698 -285927
rect 29447 -285967 30698 -285960
rect 23473 -286032 25612 -285990
rect 17406 -286184 23155 -286128
rect 22968 -286380 25227 -286367
rect 22968 -286430 23073 -286380
rect 25187 -286430 25227 -286380
rect 22968 -286498 23089 -286430
rect 25162 -286498 25227 -286430
rect 16977 -286949 17350 -286516
rect 17445 -286949 17818 -286516
rect 17913 -286949 18286 -286516
rect 18381 -286949 18754 -286516
rect 18849 -286949 19222 -286516
rect 19317 -286949 19690 -286516
rect 19785 -286949 20158 -286516
rect 20253 -286949 20626 -286516
rect 20721 -286949 21094 -286516
rect 21189 -286949 21562 -286516
rect 21657 -286949 22030 -286516
rect 22125 -286949 22604 -286516
rect 22777 -286949 22793 -286516
rect 22968 -286523 25227 -286498
rect 22361 -287110 22514 -287045
rect 16743 -289349 17116 -288916
rect 17211 -289349 17584 -288916
rect 17679 -289349 18052 -288916
rect 18147 -289349 18520 -288916
rect 18615 -289349 18988 -288916
rect 19083 -289349 19456 -288916
rect 19551 -289349 19924 -288916
rect 20019 -289349 20392 -288916
rect 20487 -289349 20860 -288916
rect 20955 -289349 21328 -288916
rect 21423 -289349 21796 -288916
rect 21891 -289349 22264 -288916
rect 22361 -289459 22409 -287110
rect 22477 -289459 22514 -287110
rect 23282 -287191 23319 -286594
rect 23500 -287191 23537 -286603
rect 23719 -287191 23756 -286592
rect 23934 -287191 23971 -286595
rect 24152 -287191 24189 -286599
rect 24374 -287191 24411 -286592
rect 24589 -287191 24626 -286595
rect 24805 -287191 24842 -286583
rect 22999 -287228 24842 -287191
rect 23584 -287339 24108 -287297
rect 22806 -287418 23307 -287402
rect 22806 -287554 22823 -287418
rect 23286 -287554 23307 -287418
rect 22806 -287570 23307 -287554
rect 22806 -288605 23007 -287570
rect 23584 -287938 23626 -287339
rect 23714 -287857 23777 -287339
rect 24065 -287428 24108 -287339
rect 24550 -287397 24592 -287228
rect 24065 -287888 24107 -287428
rect 24549 -287457 24592 -287397
rect 24176 -287514 24218 -287493
rect 24064 -287939 24107 -287888
rect 24064 -287941 24106 -287939
rect 24549 -287941 24591 -287457
rect 25570 -287654 25612 -286032
rect 26242 -286340 30542 -286311
rect 26242 -286392 26290 -286340
rect 30511 -286392 30542 -286340
rect 26242 -286419 30542 -286392
rect 30644 -286485 30698 -285967
rect 30764 -285963 30799 -285687
rect 30860 -285867 30899 -285616
rect 31201 -285767 31241 -285043
rect 31301 -285648 31341 -284710
rect 31301 -285688 33729 -285648
rect 31201 -285807 33638 -285767
rect 30860 -285906 33417 -285867
rect 30764 -285998 33285 -285963
rect 31688 -286470 32882 -286441
rect 30834 -286478 31401 -286477
rect 25699 -286864 26258 -286845
rect 25699 -286925 25723 -286864
rect 26213 -286925 26258 -286864
rect 25699 -286926 25738 -286925
rect 26202 -286926 26258 -286925
rect 25699 -286941 26258 -286926
rect 25891 -287588 25922 -287044
rect 26048 -287588 26079 -287047
rect 26437 -287588 26468 -286520
rect 26596 -287588 26627 -286511
rect 26774 -286699 26858 -286690
rect 26774 -287372 26858 -286795
rect 26774 -287481 26858 -287475
rect 26980 -287588 27011 -286519
rect 27143 -287588 27174 -286522
rect 27524 -287588 27555 -286519
rect 27682 -287588 27713 -286526
rect 28070 -287588 28101 -286510
rect 28228 -287588 28259 -286517
rect 28618 -287588 28649 -286512
rect 28768 -287588 28799 -286517
rect 29159 -286940 29190 -286518
rect 28956 -286942 29225 -286940
rect 29310 -286942 29341 -286520
rect 28956 -286971 29342 -286942
rect 28956 -287588 28987 -286971
rect 29160 -286973 29342 -286971
rect 29157 -287367 29188 -287045
rect 29216 -287360 29280 -287113
rect 29317 -287360 29348 -287041
rect 29216 -287367 29348 -287360
rect 29702 -287362 29731 -286519
rect 29862 -287362 29891 -286521
rect 30069 -286539 30698 -286485
rect 30822 -286500 31401 -286478
rect 30822 -286538 30990 -286500
rect 31307 -286531 31401 -286500
rect 31307 -286538 31346 -286531
rect 30069 -286835 30123 -286539
rect 30822 -286555 31346 -286538
rect 30822 -286769 30891 -286555
rect 30951 -286637 31203 -286602
rect 30069 -286868 30373 -286835
rect 30069 -287131 30123 -286868
rect 30951 -286913 30986 -286637
rect 30223 -286932 30986 -286913
rect 30223 -286958 31206 -286932
rect 30951 -286967 31206 -286958
rect 30309 -287074 30626 -287034
rect 30069 -287316 30173 -287131
rect 25891 -287619 28987 -287588
rect 29138 -287431 29375 -287367
rect 29138 -287588 29202 -287431
rect 29317 -287588 29348 -287431
rect 29503 -287588 29534 -287587
rect 29700 -287588 29731 -287362
rect 29861 -287588 29892 -287362
rect 29138 -287619 29892 -287588
rect 30069 -287617 30123 -287316
rect 30586 -287366 30626 -287074
rect 30309 -287404 30626 -287366
rect 30951 -287035 30986 -286967
rect 30951 -287070 31199 -287035
rect 30951 -287364 30986 -287070
rect 30951 -287399 31203 -287364
rect 30309 -287406 30605 -287404
rect 30306 -287549 30344 -287406
rect 30951 -287547 30986 -287399
rect 31325 -287471 31346 -286555
rect 31380 -287471 31401 -286531
rect 31688 -286595 31722 -286470
rect 32843 -286595 32882 -286470
rect 31688 -286651 32882 -286595
rect 31325 -287505 31401 -287471
rect 31680 -286755 31892 -286720
rect 31996 -286754 32327 -286719
rect 32426 -286754 32721 -286719
rect 31680 -286986 31715 -286755
rect 31680 -287021 31898 -286986
rect 31996 -286990 32031 -286754
rect 32426 -286987 32461 -286754
rect 31680 -287097 31715 -287021
rect 31996 -287025 32320 -286990
rect 32426 -287022 32737 -286987
rect 31996 -287093 32031 -287025
rect 32426 -287093 32461 -287022
rect 31680 -287132 31891 -287097
rect 31996 -287128 32314 -287093
rect 32426 -287128 32735 -287093
rect 31680 -287359 31715 -287132
rect 31680 -287394 31899 -287359
rect 31996 -287362 32031 -287128
rect 30951 -287582 31246 -287547
rect 30951 -287586 30986 -287582
rect 29138 -287620 29202 -287619
rect 30069 -287627 30688 -287617
rect 25570 -287696 28523 -287654
rect 30069 -287671 31157 -287627
rect 30618 -287681 31157 -287671
rect 28489 -287708 28523 -287696
rect 28489 -287742 30230 -287708
rect 30272 -287741 30443 -287708
rect 26915 -287858 30166 -287824
rect 25676 -287935 26582 -287887
rect 25676 -288393 25724 -287935
rect 26087 -287939 26571 -287935
rect 26526 -288251 26571 -287939
rect 24876 -288441 25724 -288393
rect 22659 -288635 23121 -288605
rect 22659 -288815 22690 -288635
rect 23090 -288815 23121 -288635
rect 22659 -288844 23121 -288815
rect 16345 -289604 16545 -289469
rect 22361 -289507 22514 -289459
rect 24876 -289604 24924 -288441
rect 27183 -288465 27217 -287858
rect 27402 -288455 27436 -287858
rect 27618 -288460 27652 -287858
rect 27838 -288463 27872 -287858
rect 28052 -288457 28086 -287858
rect 28272 -288452 28306 -287858
rect 28493 -288443 28527 -287858
rect 28983 -288449 29017 -287858
rect 29482 -288458 29516 -287858
rect 29707 -288456 29741 -287858
rect 29918 -288456 29952 -287858
rect 30132 -287929 30166 -287858
rect 30132 -287972 30169 -287929
rect 30135 -288456 30169 -287972
rect 30410 -288288 30443 -287741
rect 31103 -288124 31157 -287681
rect 31211 -287703 31246 -287582
rect 31211 -287738 31556 -287703
rect 31680 -287705 31715 -287394
rect 31996 -287397 32312 -287362
rect 32426 -287363 32461 -287128
rect 33250 -287363 33285 -285998
rect 31996 -287705 32031 -287397
rect 32426 -287398 33285 -287363
rect 32426 -287532 32461 -287398
rect 33378 -287530 33417 -285906
rect 32207 -287581 32461 -287532
rect 32879 -287569 33417 -287530
rect 32426 -287701 32461 -287581
rect 31211 -287947 31246 -287738
rect 31680 -287740 31893 -287705
rect 31996 -287740 32312 -287705
rect 32426 -287736 32731 -287701
rect 31680 -287947 31715 -287740
rect 31211 -287982 31558 -287947
rect 31680 -287982 31895 -287947
rect 31996 -287948 32031 -287740
rect 32426 -287944 32461 -287736
rect 31996 -287983 32310 -287948
rect 32426 -287979 32730 -287944
rect 32037 -288061 32861 -288044
rect 32037 -288116 32066 -288061
rect 32836 -288116 32861 -288061
rect 31103 -288156 31729 -288124
rect 32037 -288130 32861 -288116
rect 31124 -288157 31729 -288156
rect 31688 -288286 31729 -288157
rect 33598 -288135 33638 -285807
rect 33689 -286330 33729 -285688
rect 33689 -286370 33964 -286330
rect 33598 -288175 33936 -288135
rect 31923 -288253 33169 -288175
rect 30410 -288321 31562 -288288
rect 31124 -288529 31157 -288321
rect 31688 -288323 31990 -288286
rect 26938 -288593 30425 -288542
rect 31124 -288562 31565 -288529
rect 31594 -288568 31654 -288373
rect 31688 -288530 31729 -288323
rect 31688 -288563 31990 -288530
rect 26938 -288658 27023 -288593
rect 30391 -288658 30425 -288593
rect 26938 -288686 30425 -288658
rect 31214 -288623 32867 -288616
rect 31214 -288681 31243 -288623
rect 32843 -288681 32867 -288623
rect 31214 -288693 32867 -288681
rect 33091 -288992 33169 -288253
rect 33091 -289010 33561 -288992
rect 33091 -289229 33112 -289010
rect 33540 -289229 33561 -289010
rect 33091 -289251 33561 -289229
rect 16345 -289652 24924 -289604
rect 16345 -289669 16545 -289652
<< via1 >>
rect 29132 -282842 29402 -282710
rect 22444 -284846 22449 -283561
rect 22449 -284846 22500 -283561
rect 22500 -284846 22515 -283561
rect 22444 -285909 22449 -285345
rect 22449 -285909 22500 -285345
rect 22500 -285909 22515 -285345
rect 22444 -285914 22515 -285909
rect 22729 -283451 22966 -283158
rect 23154 -283964 25400 -283911
rect 29230 -284040 29302 -283744
rect 22740 -286051 22952 -285435
rect 23981 -285638 24303 -285574
rect 24413 -285638 25378 -285574
rect 30440 -284917 30742 -284822
rect 30857 -285527 31138 -285182
rect 23949 -285855 24451 -285798
rect 23089 -286430 25162 -286400
rect 23089 -286498 25162 -286430
rect 22604 -286949 22777 -286516
rect 22409 -287116 22477 -287110
rect 22409 -289459 22456 -287116
rect 22456 -289459 22477 -287116
rect 22823 -287554 23286 -287418
rect 26290 -286341 30511 -286340
rect 26290 -286392 30511 -286341
rect 25723 -286880 26213 -286864
rect 25723 -286925 25738 -286880
rect 25738 -286925 26202 -286880
rect 26202 -286925 26213 -286880
rect 26774 -286795 26858 -286699
rect 26774 -287475 26858 -287372
rect 31722 -286595 32843 -286470
rect 22690 -288815 23090 -288635
rect 32066 -288116 32836 -288061
rect 27023 -288658 30391 -288593
rect 31243 -288637 32843 -288623
rect 31243 -288681 32843 -288637
rect 33112 -289229 33540 -289010
<< metal2 >>
rect 38286 -282277 38605 -282252
rect 38286 -282607 38315 -282277
rect 29079 -282710 38315 -282607
rect 29079 -282842 29132 -282710
rect 29402 -282842 38315 -282710
rect 29079 -282866 38315 -282842
rect 21643 -283158 30100 -283157
rect 21643 -283450 22729 -283158
rect 21643 -283655 21936 -283450
rect 22722 -283451 22729 -283450
rect 22966 -283450 32957 -283158
rect 22966 -283451 23006 -283450
rect 29421 -283451 32957 -283450
rect 22360 -283561 22595 -283546
rect 21626 -283701 22319 -283655
rect 21626 -283951 21652 -283701
rect 22286 -283951 22319 -283701
rect 21626 -283981 22319 -283951
rect 22360 -284846 22444 -283561
rect 22515 -283849 22595 -283561
rect 29421 -283647 29988 -283451
rect 34679 -283486 36830 -283185
rect 38286 -283190 38315 -282866
rect 38576 -283190 38605 -282277
rect 38286 -283225 38605 -283190
rect 29214 -283744 29320 -283713
rect 22515 -283911 25500 -283849
rect 22515 -283964 23154 -283911
rect 25400 -283964 25500 -283911
rect 22515 -284038 25500 -283964
rect 22515 -284846 22595 -284038
rect 23187 -284504 23234 -284162
rect 23312 -284293 23386 -284038
rect 23468 -284504 23514 -284156
rect 23187 -284551 23514 -284504
rect 22360 -284861 22595 -284846
rect 23273 -284964 23358 -284828
rect 16516 -285228 23358 -284964
rect 22360 -285345 22595 -285330
rect 22360 -285914 22444 -285345
rect 22515 -285914 22595 -285345
rect 22360 -285970 22595 -285914
rect 22728 -285435 22966 -285421
rect 18233 -286032 18704 -286031
rect 22360 -286032 22515 -285970
rect 16520 -286125 16720 -286064
rect 16520 -286181 17659 -286125
rect 16520 -286264 16720 -286181
rect 18225 -286279 22515 -286032
rect 22360 -287064 22515 -286279
rect 22728 -286051 22740 -285435
rect 22952 -286051 22966 -285435
rect 23094 -285546 23358 -285228
rect 23468 -285393 23514 -284551
rect 23654 -284509 23702 -284154
rect 23776 -284301 23850 -284038
rect 23943 -284509 23988 -284144
rect 24064 -284292 24173 -284038
rect 23654 -284560 24016 -284509
rect 23620 -285546 23705 -284819
rect 23811 -285392 23862 -284560
rect 24064 -285546 24162 -284800
rect 24270 -285301 24313 -284157
rect 24384 -284289 24493 -284038
rect 24583 -284532 24626 -284158
rect 24708 -284290 24817 -284038
rect 24897 -284446 24944 -284153
rect 24504 -284552 24626 -284532
rect 24504 -284741 24522 -284552
rect 24595 -284741 24626 -284552
rect 24748 -284464 24944 -284446
rect 24748 -284653 24767 -284464
rect 24840 -284653 24944 -284464
rect 24748 -284671 24944 -284653
rect 24504 -284758 24626 -284741
rect 24386 -285546 24484 -284793
rect 24583 -285302 24626 -284758
rect 24699 -285546 24797 -284791
rect 24897 -285312 24944 -284671
rect 25029 -284490 25068 -284148
rect 25159 -284333 25251 -284038
rect 29214 -284040 29230 -283744
rect 29302 -284040 29320 -283744
rect 29421 -283860 29456 -283647
rect 29947 -283860 29988 -283647
rect 30216 -283803 31428 -283569
rect 34766 -283710 35153 -283486
rect 29421 -284012 29988 -283860
rect 25327 -284490 25374 -284155
rect 25029 -284557 25437 -284490
rect 25029 -285296 25068 -284557
rect 25141 -285546 25237 -284796
rect 25327 -285314 25374 -284557
rect 27065 -284854 27097 -284442
rect 26911 -284891 27097 -284854
rect 27366 -284452 28178 -284419
rect 27366 -285173 27399 -284452
rect 27615 -284677 27844 -284634
rect 23094 -285574 25967 -285546
rect 23094 -285638 23981 -285574
rect 24303 -285638 24413 -285574
rect 25378 -285638 25967 -285574
rect 23094 -285735 25967 -285638
rect 23066 -285799 23416 -285790
rect 23929 -285798 24465 -285788
rect 23929 -285855 23949 -285798
rect 24451 -285855 24465 -285798
rect 23929 -285869 24465 -285855
rect 23066 -285956 23416 -285939
rect 22728 -286217 22966 -286051
rect 23176 -285986 23416 -285956
rect 23176 -286126 25594 -285986
rect 22728 -286400 25356 -286217
rect 22728 -286426 23089 -286400
rect 22921 -286498 23089 -286426
rect 25162 -286498 25356 -286400
rect 22604 -286516 22777 -286508
rect 22921 -286535 25356 -286498
rect 25180 -286641 25355 -286535
rect 22992 -286816 25355 -286641
rect 22361 -287110 22514 -287064
rect 16397 -287333 16638 -287306
rect 16397 -288716 16416 -287333
rect 16602 -288716 16638 -287333
rect 21258 -288296 21935 -288273
rect 21258 -288570 21295 -288296
rect 21891 -288451 21935 -288296
rect 22361 -288451 22409 -287110
rect 21891 -288570 22409 -288451
rect 21258 -288696 22409 -288570
rect 16397 -289846 16638 -288716
rect 22361 -289459 22409 -288696
rect 22477 -288455 22514 -287110
rect 22604 -287734 22777 -286949
rect 22993 -287023 25034 -286855
rect 22993 -287402 23161 -287023
rect 22806 -287418 23516 -287402
rect 22806 -287554 22823 -287418
rect 23286 -287554 23516 -287418
rect 25180 -287438 25355 -286816
rect 22806 -287570 23516 -287554
rect 22604 -287907 23205 -287734
rect 23417 -287868 23516 -287570
rect 23032 -288201 23205 -287907
rect 23680 -288006 23787 -287539
rect 24152 -287606 24509 -287454
rect 24646 -287613 25355 -287438
rect 25454 -287675 25594 -286126
rect 25751 -286186 25967 -285735
rect 27615 -285742 27658 -284677
rect 27966 -284835 28013 -284528
rect 28145 -284713 28178 -284452
rect 28372 -284547 28478 -284517
rect 28145 -284746 28332 -284713
rect 27836 -284882 28013 -284835
rect 27836 -285662 27883 -284882
rect 28448 -284947 28478 -284547
rect 28105 -284977 28478 -284947
rect 28105 -285176 28135 -284977
rect 28325 -285814 28371 -285163
rect 28632 -285248 28676 -284482
rect 29214 -285938 29320 -284040
rect 29601 -284603 29799 -284551
rect 29601 -285815 29653 -284603
rect 30433 -284822 30742 -283803
rect 34695 -284300 35156 -284216
rect 36844 -284264 37044 -284187
rect 36758 -284363 37044 -284264
rect 36844 -284387 37044 -284363
rect 30433 -284917 30440 -284822
rect 30433 -284924 30742 -284917
rect 29760 -285582 29802 -285143
rect 30433 -286186 30741 -284924
rect 30847 -285182 31153 -285165
rect 30847 -285527 30857 -285182
rect 31138 -285365 31153 -285182
rect 34568 -285365 36846 -284986
rect 31138 -285366 36846 -285365
rect 31138 -285527 36841 -285366
rect 30847 -285535 36841 -285527
rect 33897 -285923 34233 -285535
rect 25751 -286255 30741 -286186
rect 25751 -286340 33765 -286255
rect 36830 -286315 37030 -286237
rect 25751 -286392 26290 -286340
rect 30511 -286392 33765 -286340
rect 36744 -286369 37030 -286315
rect 25751 -286470 33765 -286392
rect 36830 -286437 37030 -286369
rect 25751 -286493 31722 -286470
rect 25751 -286639 25967 -286493
rect 26303 -286632 26383 -286493
rect 25749 -286844 25967 -286639
rect 26678 -286642 26758 -286493
rect 26840 -286641 26920 -286493
rect 27227 -286649 27307 -286493
rect 27388 -286651 27468 -286493
rect 27773 -286654 27853 -286493
rect 27942 -286655 28022 -286493
rect 28317 -286655 28397 -286493
rect 28483 -286661 28563 -286493
rect 28853 -286665 28933 -286493
rect 26307 -286795 26774 -286699
rect 26858 -286795 29029 -286699
rect 29204 -286712 29308 -286493
rect 29929 -286548 29995 -286546
rect 29478 -286611 29995 -286548
rect 29478 -286741 29541 -286611
rect 25749 -286846 28906 -286844
rect 25705 -286864 28906 -286846
rect 25705 -286925 25723 -286864
rect 26213 -286925 28906 -286864
rect 25705 -286943 28906 -286925
rect 25749 -287062 28906 -286943
rect 28948 -286905 29029 -286795
rect 29064 -286804 29541 -286741
rect 29601 -286797 29667 -286611
rect 29759 -286835 29825 -286659
rect 29929 -286788 29995 -286611
rect 30110 -286595 31722 -286493
rect 32843 -286595 33765 -286470
rect 30110 -286620 33765 -286595
rect 30110 -286786 30207 -286620
rect 29759 -286901 30135 -286835
rect 28948 -286907 29044 -286905
rect 28948 -287003 29476 -286907
rect 25752 -287203 25862 -287062
rect 25937 -287372 26047 -287154
rect 26124 -287216 26234 -287062
rect 26293 -287223 26403 -287062
rect 26482 -287372 26592 -287170
rect 26658 -287238 26768 -287062
rect 26870 -287292 26961 -287062
rect 25937 -287475 26774 -287372
rect 26858 -287475 26865 -287372
rect 27024 -287373 27125 -287120
rect 27185 -287296 27276 -287062
rect 27418 -287291 27511 -287062
rect 27584 -287373 27677 -287119
rect 27737 -287300 27830 -287062
rect 27957 -287286 28050 -287062
rect 28112 -287373 28205 -287128
rect 28287 -287291 28380 -287062
rect 28498 -287291 28591 -287062
rect 28663 -287373 28756 -287128
rect 28835 -287282 28906 -287062
rect 29042 -287288 29138 -287003
rect 29380 -287303 29476 -287003
rect 29587 -287060 30003 -286969
rect 29587 -287373 29678 -287060
rect 27024 -287466 29678 -287373
rect 29747 -287363 29838 -287166
rect 29912 -287318 30003 -287060
rect 30059 -287039 30135 -286901
rect 30273 -286965 30334 -286659
rect 30393 -286784 30490 -286620
rect 30059 -287115 30551 -287039
rect 30483 -287244 30551 -287115
rect 30147 -287326 30451 -287265
rect 30826 -287363 30888 -286761
rect 31051 -287363 31097 -286751
rect 29747 -287455 31097 -287363
rect 29747 -287456 31079 -287455
rect 27034 -287471 29678 -287466
rect 29123 -287554 29212 -287553
rect 23935 -287827 27068 -287675
rect 23938 -287923 24374 -287827
rect 23680 -288164 24921 -288006
rect 25066 -288164 26453 -288006
rect 23680 -288167 23787 -288164
rect 26639 -288201 26731 -287972
rect 26916 -287990 27068 -287827
rect 28678 -287680 28827 -287611
rect 28678 -287890 28703 -287680
rect 28807 -287890 28827 -287680
rect 28678 -287913 28827 -287890
rect 29123 -287639 29409 -287554
rect 26916 -288148 28651 -287990
rect 27044 -288149 28651 -288148
rect 23032 -288374 26731 -288201
rect 26639 -288377 26731 -288374
rect 23847 -288455 24070 -288450
rect 27270 -288455 27366 -288209
rect 27698 -288455 27794 -288202
rect 28137 -288455 28233 -288201
rect 28566 -288455 28662 -288201
rect 28812 -288455 28895 -287992
rect 29123 -288388 29212 -287639
rect 30306 -287752 30352 -287522
rect 29342 -288187 30347 -288017
rect 30980 -288128 31034 -287534
rect 31224 -287538 31272 -286746
rect 31746 -287301 31816 -286620
rect 31768 -287306 31816 -287301
rect 31224 -287586 31543 -287538
rect 31269 -287942 31330 -287788
rect 31442 -287822 31490 -287586
rect 31884 -287615 31932 -286810
rect 32071 -287308 32140 -286620
rect 32071 -287309 32135 -287308
rect 32204 -287532 32252 -286807
rect 32311 -287308 32388 -286620
rect 32471 -287301 32545 -286620
rect 32324 -287313 32388 -287308
rect 32497 -287309 32545 -287301
rect 32623 -287526 32671 -286806
rect 32730 -287311 32812 -286620
rect 33427 -287044 33765 -286620
rect 33886 -287044 34050 -286958
rect 33427 -287073 34050 -287044
rect 33427 -287362 33758 -287073
rect 33974 -287362 34050 -287073
rect 33427 -287392 34050 -287362
rect 33886 -287524 34050 -287392
rect 32204 -287581 32457 -287532
rect 32623 -287580 32887 -287526
rect 31884 -287663 31964 -287615
rect 31599 -287942 31794 -287770
rect 31916 -287889 31964 -287663
rect 32036 -287942 32116 -287786
rect 32204 -287799 32252 -287581
rect 32340 -287942 32543 -287783
rect 32623 -287801 32671 -287580
rect 32757 -287942 32820 -287780
rect 31181 -288061 32918 -287942
rect 31181 -288098 32066 -288061
rect 32024 -288116 32066 -288098
rect 32836 -288116 32918 -288061
rect 36815 -288112 37015 -288045
rect 30980 -288182 31958 -288128
rect 32024 -288138 32918 -288116
rect 30295 -288210 30347 -288187
rect 29554 -288455 29660 -288227
rect 29996 -288455 30102 -288236
rect 30295 -288256 31807 -288210
rect 31436 -288344 31713 -288290
rect 31276 -288455 31340 -288369
rect 22477 -289258 22515 -288455
rect 23293 -288472 31340 -288455
rect 22659 -288635 23121 -288606
rect 22659 -288815 22690 -288635
rect 23090 -288815 23121 -288635
rect 23293 -288679 25084 -288472
rect 25590 -288533 31340 -288472
rect 31436 -288493 31520 -288344
rect 31594 -288533 31675 -288389
rect 25590 -288577 31675 -288533
rect 31751 -288527 31807 -288256
rect 31904 -288495 31958 -288182
rect 32299 -288143 32916 -288138
rect 32299 -288337 32413 -288143
rect 32786 -288337 32916 -288143
rect 36711 -288173 37015 -288112
rect 36815 -288245 37015 -288173
rect 37660 -288114 38614 -288081
rect 32067 -288527 32123 -288356
rect 25590 -288593 31674 -288577
rect 31751 -288583 32123 -288527
rect 32299 -288550 32916 -288337
rect 37660 -288362 37705 -288114
rect 38569 -288362 38614 -288114
rect 37660 -288400 38614 -288362
rect 25590 -288658 27023 -288593
rect 30391 -288612 31674 -288593
rect 32299 -288612 33906 -288550
rect 30391 -288623 33906 -288612
rect 30391 -288658 31243 -288623
rect 25590 -288679 31243 -288658
rect 23293 -288681 31243 -288679
rect 32843 -288681 33906 -288623
rect 23293 -288696 33906 -288681
rect 23293 -288697 32880 -288696
rect 23293 -288698 31674 -288697
rect 22659 -288844 23121 -288815
rect 23294 -289258 23836 -288698
rect 37676 -288778 37759 -288400
rect 28637 -288790 37759 -288778
rect 28637 -288849 28651 -288790
rect 28898 -288849 37759 -288790
rect 28637 -288861 37759 -288849
rect 38283 -288802 38605 -288781
rect 38283 -288992 38309 -288802
rect 33089 -289010 38309 -288992
rect 33089 -289229 33112 -289010
rect 33540 -289229 38309 -289010
rect 33089 -289251 38309 -289229
rect 22477 -289459 23836 -289258
rect 22361 -289846 23836 -289459
rect 38283 -289668 38309 -289251
rect 38582 -289668 38605 -288802
rect 38283 -289695 38605 -289668
rect 16282 -290388 23836 -289846
rect 16289 -290641 16831 -290388
rect 1322 -290642 16831 -290641
rect 1313 -290662 16831 -290642
rect 1313 -291165 1338 -290662
rect 1610 -291165 16831 -290662
rect 1313 -291183 16831 -291165
rect 1313 -291185 1631 -291183
<< via2 >>
rect 21652 -283951 22286 -283701
rect 38315 -283190 38576 -282277
rect 24522 -284741 24595 -284552
rect 24767 -284653 24840 -284464
rect 29456 -283860 29947 -283647
rect 23066 -285939 23416 -285799
rect 23949 -285855 24451 -285798
rect 16416 -288716 16602 -287333
rect 21295 -288570 21891 -288296
rect 24921 -288164 25066 -288006
rect 28703 -287890 28807 -287680
rect 33758 -287362 33974 -287073
rect 22690 -288815 23090 -288635
rect 25084 -288679 25590 -288472
rect 37705 -288362 38569 -288114
rect 28651 -288849 28898 -288790
rect 38309 -289668 38582 -288802
rect 1338 -291165 1610 -290662
<< metal3 >>
rect 38286 -282277 38605 -282252
rect 38286 -283190 38315 -282277
rect 38576 -283190 38605 -282277
rect 38286 -283225 38605 -283190
rect 24750 -283541 25100 -283526
rect 24750 -283617 24767 -283541
rect 25081 -283617 25100 -283541
rect 24750 -283631 25100 -283617
rect 21626 -283701 22386 -283669
rect 21626 -283951 21652 -283701
rect 22286 -283951 22386 -283701
rect 21626 -283981 22386 -283951
rect 24750 -284447 24811 -283631
rect 28953 -283647 29989 -283631
rect 24920 -283728 25370 -283705
rect 24749 -284464 24860 -284447
rect 24504 -284552 24615 -284532
rect 24504 -284741 24522 -284552
rect 24595 -284741 24615 -284552
rect 24749 -284653 24767 -284464
rect 24840 -284653 24860 -284464
rect 24920 -284604 25068 -283728
rect 25317 -284604 25370 -283728
rect 24920 -284627 25370 -284604
rect 28953 -283860 29456 -283647
rect 29947 -283860 29989 -283647
rect 28953 -283897 29989 -283860
rect 24749 -284674 24860 -284653
rect 24504 -284759 24615 -284741
rect 24508 -285582 24576 -284759
rect 24508 -285595 24803 -285582
rect 24508 -285694 24576 -285595
rect 24790 -285694 24803 -285595
rect 22189 -285723 22809 -285701
rect 24508 -285707 24803 -285694
rect 16394 -285961 17240 -285925
rect 16394 -286321 16440 -285961
rect 17201 -286321 17240 -285961
rect 22189 -285999 22225 -285723
rect 22783 -285799 22809 -285723
rect 23061 -285799 23421 -285794
rect 22783 -285939 23066 -285799
rect 23416 -285939 23421 -285799
rect 23929 -285798 24465 -285788
rect 23929 -285855 23949 -285798
rect 24451 -285827 24465 -285798
rect 24540 -285827 24863 -285801
rect 24451 -285829 24863 -285827
rect 24451 -285855 24568 -285829
rect 23929 -285869 24568 -285855
rect 22783 -285999 22809 -285939
rect 23061 -285944 23421 -285939
rect 23930 -285971 24568 -285869
rect 22189 -286022 22809 -285999
rect 18233 -286278 18704 -286031
rect 24540 -286134 24568 -285971
rect 24832 -286134 24863 -285829
rect 24540 -286158 24863 -286134
rect 16394 -286357 17240 -286321
rect 16397 -287333 16637 -286357
rect 16397 -288716 16416 -287333
rect 16602 -288716 16637 -287333
rect 24923 -287994 25068 -284627
rect 25248 -284977 25464 -284974
rect 25179 -285016 25501 -284977
rect 25179 -285880 25218 -285016
rect 25463 -285880 25501 -285016
rect 28953 -285522 29219 -283897
rect 25179 -285917 25501 -285880
rect 28899 -285564 29219 -285522
rect 25217 -286281 25464 -285917
rect 25183 -286323 25488 -286281
rect 25183 -287128 25224 -286323
rect 25445 -287128 25488 -286323
rect 28899 -286699 28949 -285564
rect 29174 -286699 29219 -285564
rect 28899 -286745 29219 -286699
rect 33956 -286411 34284 -286385
rect 33956 -287044 33985 -286411
rect 25183 -287175 25488 -287128
rect 33725 -287073 33985 -287044
rect 24913 -288006 25074 -287994
rect 24913 -288164 24921 -288006
rect 25066 -288164 25074 -288006
rect 24913 -288177 25074 -288164
rect 21258 -288296 22022 -288274
rect 21258 -288570 21295 -288296
rect 21891 -288303 22022 -288296
rect 21899 -288568 22022 -288303
rect 25217 -288454 25464 -287175
rect 33725 -287362 33758 -287073
rect 33974 -287362 33985 -287073
rect 33725 -287391 33985 -287362
rect 28679 -287680 28829 -287661
rect 28679 -287890 28703 -287680
rect 28807 -287890 28829 -287680
rect 33956 -287739 33985 -287391
rect 34247 -287739 34284 -286411
rect 33956 -287771 34284 -287739
rect 21891 -288570 22022 -288568
rect 21258 -288600 22022 -288570
rect 25059 -288472 25615 -288454
rect 16397 -288754 16637 -288716
rect 22659 -288627 23121 -288605
rect 22659 -288810 22684 -288627
rect 23094 -288810 23121 -288627
rect 25059 -288679 25084 -288472
rect 25590 -288679 25615 -288472
rect 25059 -288699 25615 -288679
rect 28679 -288778 28829 -287890
rect 37660 -288114 38614 -288081
rect 37660 -288362 37705 -288114
rect 38569 -288362 38614 -288114
rect 37660 -288400 38614 -288362
rect 22659 -288815 22690 -288810
rect 23090 -288815 23121 -288810
rect 22659 -288844 23121 -288815
rect 28637 -288790 28914 -288778
rect 28637 -288849 28651 -288790
rect 28898 -288849 28914 -288790
rect 28637 -288861 28914 -288849
rect 38283 -288802 38605 -288781
rect 38283 -289668 38309 -288802
rect 38582 -289668 38605 -288802
rect 38283 -289695 38605 -289668
rect 1313 -290662 1631 -290642
rect 1313 -291165 1338 -290662
rect 1610 -291165 1631 -290662
rect 1313 -291185 1631 -291165
<< via3 >>
rect 38315 -283190 38576 -282277
rect 24767 -283617 25081 -283541
rect 21652 -283951 22286 -283701
rect 25068 -284604 25317 -283728
rect 24576 -285694 24790 -285595
rect 16440 -286321 17201 -285961
rect 22225 -285999 22783 -285723
rect 24568 -286134 24832 -285829
rect 25218 -285880 25463 -285016
rect 25224 -287128 25445 -286323
rect 28949 -286699 29174 -285564
rect 21300 -288568 21891 -288303
rect 21891 -288568 21899 -288303
rect 33985 -287739 34247 -286411
rect 22684 -288635 23094 -288627
rect 22684 -288810 22690 -288635
rect 22690 -288810 23090 -288635
rect 23090 -288810 23094 -288635
rect 37705 -288362 38569 -288114
rect 38309 -289668 38582 -288802
rect 1338 -291165 1610 -290662
<< metal4 >>
rect 38284 -276864 38606 -276836
rect 38284 -277025 38312 -276864
rect 37750 -277347 38312 -277025
rect 38284 -277490 38312 -277347
rect 38575 -277490 38606 -276864
rect 38284 -277532 38606 -277490
rect 1315 -278744 1635 -278710
rect 1315 -279007 1340 -278744
rect 1312 -279111 1340 -279007
rect 1315 -279302 1340 -279111
rect 1600 -278999 1635 -278744
rect 1600 -279103 2168 -278999
rect 1600 -279302 1635 -279103
rect 1315 -279342 1635 -279302
rect 38282 -281174 38604 -281146
rect 38282 -281323 38310 -281174
rect 37750 -281645 38310 -281323
rect 38282 -281800 38310 -281645
rect 38573 -281323 38604 -281174
rect 38573 -281645 38606 -281323
rect 38573 -281800 38604 -281645
rect 38282 -281841 38604 -281800
rect 38286 -282277 38605 -282252
rect 1315 -283060 1635 -283026
rect 1315 -283319 1340 -283060
rect 1313 -283423 1340 -283319
rect 1315 -283618 1340 -283423
rect 1600 -283311 1635 -283060
rect 38286 -283190 38315 -282277
rect 38576 -283190 38605 -282277
rect 38286 -283225 38605 -283190
rect 1600 -283415 2154 -283311
rect 1600 -283618 1635 -283415
rect 1315 -283658 1635 -283618
rect 24749 -283541 29224 -283527
rect 24749 -283617 24767 -283541
rect 25081 -283617 29224 -283541
rect 24749 -283631 29224 -283617
rect 21626 -283687 22389 -283654
rect 21626 -283701 21692 -283687
rect 21626 -283951 21652 -283701
rect 22345 -283936 22389 -283687
rect 28903 -283700 29224 -283631
rect 22286 -283951 22389 -283936
rect 21626 -283983 22389 -283951
rect 25038 -283728 25505 -283705
rect 25038 -284604 25068 -283728
rect 25317 -283745 25505 -283728
rect 25475 -284574 25505 -283745
rect 25317 -284604 25505 -284574
rect 25038 -284626 25505 -284604
rect 28903 -283745 29223 -283700
rect 28903 -284608 28946 -283745
rect 29183 -284608 29223 -283745
rect 25038 -284627 25488 -284626
rect 28903 -284649 29223 -284608
rect 25179 -285012 25499 -284973
rect 24528 -285595 25097 -285583
rect 24528 -285694 24576 -285595
rect 24790 -285694 25097 -285595
rect 22189 -285723 22809 -285701
rect 24528 -285707 25097 -285694
rect 16396 -285961 17682 -285926
rect 16396 -286321 16440 -285961
rect 17201 -286321 17682 -285961
rect 22189 -285999 22225 -285723
rect 22783 -285999 22809 -285723
rect 22189 -286022 22809 -285999
rect 24542 -285828 24862 -285801
rect 24542 -286135 24568 -285828
rect 24834 -286135 24862 -285828
rect 24973 -285992 25097 -285707
rect 25179 -285876 25217 -285012
rect 25458 -285016 25499 -285012
rect 25463 -285603 25499 -285016
rect 28897 -285563 29217 -285524
rect 25179 -285880 25218 -285876
rect 25463 -285880 25710 -285603
rect 25179 -285922 25710 -285880
rect 25430 -285925 25710 -285922
rect 24973 -286116 28757 -285992
rect 24542 -286162 24862 -286135
rect 25465 -286278 25668 -286275
rect 16396 -286362 17682 -286321
rect 25185 -286323 25668 -286278
rect 25185 -286328 25224 -286323
rect 25445 -286328 25668 -286323
rect 25185 -287129 25223 -286328
rect 25464 -286593 25668 -286328
rect 25464 -287129 25505 -286593
rect 25185 -287178 25505 -287129
rect 25183 -287584 25503 -287543
rect 21258 -288303 22021 -288273
rect 21258 -288318 21300 -288303
rect 21899 -288318 22021 -288303
rect 21258 -288556 21295 -288318
rect 21969 -288556 22021 -288318
rect 25183 -288385 25227 -287584
rect 25468 -288385 25503 -287584
rect 28633 -287544 28757 -286116
rect 28897 -286713 28932 -285563
rect 29182 -285912 29217 -285563
rect 29182 -286228 29472 -285912
rect 29182 -286713 29217 -286228
rect 28897 -286749 29217 -286713
rect 33957 -286394 34277 -286387
rect 33957 -286411 34435 -286394
rect 33957 -286445 33985 -286411
rect 28893 -287544 29213 -287541
rect 28633 -287583 29213 -287544
rect 28633 -287668 28941 -287583
rect 25183 -288425 25503 -288385
rect 28893 -288453 28941 -287668
rect 29177 -288453 29213 -287583
rect 33957 -287727 33982 -286445
rect 34247 -286719 34435 -286411
rect 33957 -287739 33985 -287727
rect 34247 -287739 34277 -286719
rect 33957 -287783 34277 -287739
rect 28893 -288490 29213 -288453
rect 33308 -287977 33629 -287947
rect 21258 -288568 21300 -288556
rect 21899 -288568 22021 -288556
rect 21258 -288602 22021 -288568
rect 22659 -288598 23121 -288596
rect 22658 -288627 23121 -288598
rect 1313 -288702 1633 -288668
rect 1313 -288965 1338 -288702
rect 1312 -289069 1338 -288965
rect 1313 -289260 1338 -289069
rect 1598 -288941 1633 -288702
rect 22658 -288810 22684 -288627
rect 23094 -288716 23121 -288627
rect 33308 -288700 33332 -287977
rect 33605 -288700 33629 -287977
rect 37659 -288114 38612 -288081
rect 37659 -288119 37705 -288114
rect 37659 -288361 37704 -288119
rect 37659 -288362 37705 -288361
rect 38569 -288362 38612 -288114
rect 37659 -288401 38612 -288362
rect 33308 -288716 33629 -288700
rect 23094 -288810 33629 -288716
rect 22658 -288841 33629 -288810
rect 23094 -288846 33629 -288841
rect 38283 -288802 38605 -288781
rect 1598 -289045 2115 -288941
rect 1598 -289260 1633 -289045
rect 1313 -289300 1633 -289260
rect 38283 -289668 38309 -288802
rect 38582 -289668 38605 -288802
rect 38283 -289695 38605 -289668
rect 38278 -290587 38600 -290559
rect 1313 -290662 1631 -290642
rect 1313 -291165 1338 -290662
rect 1610 -291165 1631 -290662
rect 38278 -290729 38306 -290587
rect 37747 -291051 38306 -290729
rect 1313 -291185 1631 -291165
rect 38278 -291213 38306 -291051
rect 38569 -290729 38600 -290587
rect 38569 -291051 38603 -290729
rect 38569 -291213 38600 -291051
rect 38278 -291254 38600 -291213
rect 1312 -293050 1633 -293016
rect 1312 -293277 1337 -293050
rect 1311 -293381 1337 -293277
rect 1312 -293608 1337 -293381
rect 1597 -293253 1633 -293050
rect 1597 -293357 2114 -293253
rect 1597 -293608 1633 -293357
rect 1312 -293648 1633 -293608
rect 38282 -294857 38604 -294829
rect 38282 -295022 38310 -294857
rect 37749 -295344 38310 -295022
rect 38282 -295483 38310 -295344
rect 38573 -295022 38604 -294857
rect 38573 -295344 38605 -295022
rect 38573 -295483 38604 -295344
rect 38282 -295524 38604 -295483
<< via4 >>
rect 38312 -277490 38575 -276864
rect 1340 -279302 1600 -278744
rect 38310 -281800 38573 -281174
rect 1340 -283618 1600 -283060
rect 38315 -283190 38576 -282277
rect 21692 -283701 22345 -283687
rect 21692 -283936 22286 -283701
rect 22286 -283936 22345 -283701
rect 25237 -284574 25317 -283745
rect 25317 -284574 25475 -283745
rect 28946 -284608 29183 -283745
rect 16440 -286321 17201 -285961
rect 22225 -285996 22783 -285725
rect 24568 -285829 24834 -285828
rect 24568 -286134 24832 -285829
rect 24832 -286134 24834 -285829
rect 24568 -286135 24834 -286134
rect 25217 -285016 25458 -285012
rect 25217 -285876 25218 -285016
rect 25218 -285876 25458 -285016
rect 25223 -287128 25224 -286328
rect 25224 -287128 25445 -286328
rect 25445 -287128 25464 -286328
rect 25223 -287129 25464 -287128
rect 21295 -288556 21300 -288318
rect 21300 -288556 21899 -288318
rect 21899 -288556 21969 -288318
rect 25227 -288385 25468 -287584
rect 28932 -285564 29182 -285563
rect 28932 -286699 28949 -285564
rect 28949 -286699 29174 -285564
rect 29174 -286699 29182 -285564
rect 28932 -286713 29182 -286699
rect 28941 -288453 29177 -287583
rect 33982 -287727 33985 -286445
rect 33985 -287727 34225 -286445
rect 1338 -289260 1598 -288702
rect 33332 -288700 33605 -287977
rect 37704 -288361 37705 -288119
rect 37705 -288361 38568 -288119
rect 38309 -289668 38582 -288802
rect 1338 -291165 1610 -290662
rect 38306 -291213 38569 -290587
rect 1337 -293608 1597 -293050
rect 38310 -295483 38573 -294857
<< metal5 >>
rect 38285 -274945 38605 -274935
rect 37932 -275265 38605 -274945
rect 38285 -276836 38605 -275265
rect 38284 -276864 38606 -276836
rect 1312 -277345 1967 -277025
rect 1312 -278710 1632 -277345
rect 38284 -277490 38312 -276864
rect 38575 -277490 38606 -276864
rect 38284 -277532 38606 -277490
rect 1312 -278744 1635 -278710
rect 1312 -279302 1340 -278744
rect 1600 -279302 1635 -278744
rect 38285 -279243 38605 -277532
rect 1312 -279342 1635 -279302
rect 1312 -281323 1632 -279342
rect 37916 -279563 38605 -279243
rect 38285 -281145 38605 -279563
rect 38283 -281146 38605 -281145
rect 38282 -281174 38605 -281146
rect 1312 -281643 1975 -281323
rect 1312 -283026 1632 -281643
rect 38282 -281800 38310 -281174
rect 38573 -281800 38605 -281174
rect 38282 -281841 38605 -281800
rect 38285 -282277 38605 -281841
rect 1312 -283060 1635 -283026
rect 1312 -283618 1340 -283060
rect 1600 -283618 1635 -283060
rect 38285 -283190 38315 -282277
rect 38576 -283190 38605 -282277
rect 38285 -283254 38605 -283190
rect 1312 -283658 1635 -283618
rect 1312 -288668 1632 -283658
rect 21636 -283687 23227 -283658
rect 21636 -283936 21692 -283687
rect 22345 -283936 23227 -283687
rect 21636 -283978 23227 -283936
rect 25185 -283745 25505 -283705
rect 25185 -284287 25237 -283745
rect 24782 -284574 25237 -284287
rect 25475 -284574 25505 -283745
rect 28903 -283745 29223 -283700
rect 28903 -284329 28946 -283745
rect 24782 -284607 25505 -284574
rect 25185 -284626 25505 -284607
rect 28462 -284608 28946 -284329
rect 29183 -284608 29223 -283745
rect 28462 -284649 29223 -284608
rect 25183 -285012 25503 -284973
rect 21665 -285725 22809 -285701
rect 16396 -285927 17220 -285926
rect 16396 -285961 18116 -285927
rect 16396 -286321 16440 -285961
rect 17201 -286321 18116 -285961
rect 21665 -285996 22225 -285725
rect 22783 -285996 22809 -285725
rect 21665 -286022 22809 -285996
rect 24542 -285828 24862 -285803
rect 24542 -286135 24568 -285828
rect 24834 -286135 24862 -285828
rect 25183 -285876 25217 -285012
rect 25458 -285602 25503 -285012
rect 28897 -285563 29217 -285524
rect 25458 -285876 26311 -285602
rect 25183 -285922 26311 -285876
rect 24542 -286257 24862 -286135
rect 16396 -286362 18116 -286321
rect 25185 -286328 26349 -286278
rect 25185 -287129 25223 -286328
rect 25464 -286598 26349 -286328
rect 25464 -287129 25505 -286598
rect 28897 -286713 28932 -285563
rect 29182 -285911 29217 -285563
rect 29182 -286231 29914 -285911
rect 29182 -286713 29219 -286231
rect 28897 -286749 29219 -286713
rect 33957 -286445 35027 -286387
rect 25185 -287178 25505 -287129
rect 24721 -287584 25503 -287543
rect 24721 -287863 25227 -287584
rect 21258 -288318 22908 -288280
rect 21258 -288556 21295 -288318
rect 21969 -288556 22908 -288318
rect 25183 -288385 25227 -287863
rect 25468 -288385 25503 -287584
rect 28385 -287583 29213 -287541
rect 28385 -287861 28941 -287583
rect 25183 -288425 25503 -288385
rect 28893 -288453 28941 -287861
rect 29177 -288453 29213 -287583
rect 33957 -287727 33982 -286445
rect 34225 -286707 35027 -286445
rect 34225 -287727 34277 -286707
rect 28893 -288490 29213 -288453
rect 33308 -287943 33628 -287777
rect 33957 -287783 34277 -287727
rect 33308 -287977 33631 -287943
rect 21258 -288600 22908 -288556
rect 1312 -288702 1633 -288668
rect 1312 -289260 1338 -288702
rect 1598 -289260 1633 -288702
rect 33308 -288700 33332 -287977
rect 33605 -288700 33631 -287977
rect 38292 -288081 38612 -287643
rect 37659 -288119 38612 -288081
rect 37659 -288361 37704 -288119
rect 38568 -288361 38612 -288119
rect 37659 -288401 38612 -288361
rect 33308 -288728 33631 -288700
rect 38285 -288777 38605 -288730
rect 38285 -288781 38607 -288777
rect 1312 -289300 1633 -289260
rect 38283 -288802 38607 -288781
rect 1312 -290634 1632 -289300
rect 38283 -289668 38309 -288802
rect 38582 -289668 38607 -288802
rect 38283 -289695 38607 -289668
rect 38285 -289700 38607 -289695
rect 38285 -290558 38605 -289700
rect 38279 -290559 38605 -290558
rect 38278 -290587 38605 -290559
rect 1312 -290662 1636 -290634
rect 1312 -291165 1338 -290662
rect 1610 -290727 1636 -290662
rect 1610 -291047 1971 -290727
rect 1610 -291165 1636 -291047
rect 1312 -291188 1636 -291165
rect 1312 -293050 1632 -291188
rect 38278 -291213 38306 -290587
rect 38569 -291213 38605 -290587
rect 38278 -291254 38605 -291213
rect 38285 -292807 38605 -291254
rect 1312 -293608 1337 -293050
rect 1597 -293608 1632 -293050
rect 37916 -293127 38605 -292807
rect 1312 -295025 1632 -293608
rect 38285 -294828 38605 -293127
rect 38283 -294829 38605 -294828
rect 38282 -294857 38605 -294829
rect 1312 -295345 1980 -295025
rect 38282 -295483 38310 -294857
rect 38573 -295483 38605 -294857
rect 38282 -295524 38605 -295483
rect 38285 -297105 38605 -295524
rect 37916 -297425 38605 -297105
rect 38285 -297437 38605 -297425
<< comment >>
rect 24359 -284563 24362 -284505
rect 24280 -284564 24362 -284563
use por_output_buffer  por_output_buffer_0
timestamp 1717613630
transform 1 0 549 0 -1 -572311
box 33352 -286528 36282 -285202
use por_output_buffer  por_output_buffer_1
timestamp 1717613630
transform 1 0 534 0 1 -2177
box 33352 -286528 36282 -285202
use por_output_driver_h  por_output_driver_h_0
timestamp 1717613630
transform 1 0 8288 0 1 7808
box 26862 -292924 28562 -291020
use por_via_2cut  por_via_2cut_0
timestamp 1717613630
transform 0 1 40548 -1 0 -271091
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_1
timestamp 1717613630
transform 0 1 34819 -1 0 -271057
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_2
timestamp 1717613630
transform 0 1 39669 -1 0 -271684
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_3
timestamp 1717613630
transform 0 1 40452 -1 0 -271090
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_4
timestamp 1717613630
transform 0 1 40228 -1 0 -271089
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_5
timestamp 1717613630
transform 0 1 40129 -1 0 -271089
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_6
timestamp 1717613630
transform 0 1 40030 -1 0 -271090
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_7
timestamp 1717613630
transform 0 1 39813 -1 0 -271092
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_8
timestamp 1717613630
transform 0 1 39715 -1 0 -271092
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_9
timestamp 1717613630
transform 0 1 39135 -1 0 -271087
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_10
timestamp 1717613630
transform 0 1 38077 -1 0 -271094
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_11
timestamp 1717613630
transform 0 1 37860 -1 0 -271087
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_12
timestamp 1717613630
transform 0 1 37700 -1 0 -271090
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_13
timestamp 1717613630
transform 0 1 39016 -1 0 -270657
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_14
timestamp 1717613630
transform 0 1 40645 -1 0 -270711
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_15
timestamp 1717613630
transform 0 1 40547 -1 0 -270710
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_16
timestamp 1717613630
transform 0 1 40450 -1 0 -270714
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_17
timestamp 1717613630
transform 0 1 40227 -1 0 -270713
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_18
timestamp 1717613630
transform 0 1 40130 -1 0 -270711
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_19
timestamp 1717613630
transform 0 1 40035 -1 0 -270714
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_20
timestamp 1717613630
transform 0 1 39807 -1 0 -270710
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_21
timestamp 1717613630
transform 0 1 39713 -1 0 -270711
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_22
timestamp 1717613630
transform 0 1 39123 -1 0 -270653
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_23
timestamp 1717613630
transform 0 1 40644 -1 0 -271091
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_24
timestamp 1717613630
transform 0 1 40543 -1 0 -271688
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_25
timestamp 1717613630
transform 0 1 39842 -1 0 -271683
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_26
timestamp 1717613630
transform -1 0 47817 0 -1 -296219
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_27
timestamp 1717613630
transform 0 1 40234 -1 0 -271686
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_28
timestamp 1717613630
transform 0 1 39987 -1 0 -271689
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_29
timestamp 1717613630
transform 0 1 40119 -1 0 -271686
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_30
timestamp 1717613630
transform 0 1 39526 -1 0 -271690
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_31
timestamp 1717613630
transform 0 1 39367 -1 0 -271686
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_32
timestamp 1717613630
transform 0 1 37941 -1 0 -272153
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_33
timestamp 1717613630
transform 0 1 40419 -1 0 -271689
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_34
timestamp 1717613630
transform 0 1 40683 -1 0 -271691
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_35
timestamp 1717613630
transform 0 1 39994 -1 0 -272266
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_36
timestamp 1717613630
transform 0 1 39834 -1 0 -272274
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_37
timestamp 1717613630
transform 0 1 39683 -1 0 -272266
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_38
timestamp 1717613630
transform 0 1 39527 -1 0 -272297
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_39
timestamp 1717613630
transform 0 1 39370 -1 0 -272272
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_40
timestamp 1717613630
transform 0 1 37535 -1 0 -271088
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_41
timestamp 1717613630
transform 0 1 37321 -1 0 -271061
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_42
timestamp 1717613630
transform 0 1 36990 -1 0 -270565
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_43
timestamp 1717613630
transform 0 1 36989 -1 0 -271052
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_44
timestamp 1717613630
transform 0 1 36774 -1 0 -271052
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_45
timestamp 1717613630
transform 0 1 36612 -1 0 -271054
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_46
timestamp 1717613630
transform 0 1 36455 -1 0 -271049
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_47
timestamp 1717613630
transform 0 1 36225 -1 0 -271059
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_48
timestamp 1717613630
transform 0 1 36067 -1 0 -271059
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_49
timestamp 1717613630
transform 0 1 35906 -1 0 -271050
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_50
timestamp 1717613630
transform 0 1 35133 -1 0 -271055
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_51
timestamp 1717613630
transform 0 1 34980 -1 0 -271061
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_52
timestamp 1717613630
transform 0 1 39008 -1 0 -271090
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_53
timestamp 1717613630
transform 0 1 38331 -1 0 -270571
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_54
timestamp 1717613630
transform 0 1 38203 -1 0 -270565
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_55
timestamp 1717613630
transform 0 1 37540 -1 0 -270577
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_56
timestamp 1717613630
transform 0 1 38418 -1 0 -271024
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_57
timestamp 1717613630
transform 0 1 38320 -1 0 -271091
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_58
timestamp 1717613630
transform 0 1 39207 -1 0 -272279
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_59
timestamp 1717613630
transform 0 1 38169 -1 0 -271945
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_60
timestamp 1717613630
transform 0 1 37733 -1 0 -271949
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_61
timestamp 1717613630
transform 0 1 37287 -1 0 -271951
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_62
timestamp 1717613630
transform 0 1 35216 -1 0 -272142
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_63
timestamp 1717613630
transform 0 1 38080 -1 0 -270555
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_64
timestamp 1717613630
transform 0 1 37691 -1 0 -270562
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_65
timestamp 1717613630
transform 0 1 37861 -1 0 -270567
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_66
timestamp 1717613630
transform 0 1 39206 -1 0 -271694
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_67
timestamp 1717613630
transform 0 1 32106 -1 0 -271386
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_68
timestamp 1717613630
transform 0 1 32589 -1 0 -271376
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_69
timestamp 1717613630
transform 0 1 37149 -1 0 -270490
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_70
timestamp 1717613630
transform 0 1 37311 -1 0 -270568
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_71
timestamp 1717613630
transform 0 1 35526 -1 0 -271063
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_72
timestamp 1717613630
transform 0 1 35687 -1 0 -271059
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_73
timestamp 1717613630
transform 0 1 35359 -1 0 -271059
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_74
timestamp 1717613630
transform 0 1 36607 -1 0 -270567
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_75
timestamp 1717613630
transform 0 1 36064 -1 0 -270567
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_76
timestamp 1717613630
transform 0 1 35521 -1 0 -270567
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_77
timestamp 1717613630
transform 0 1 34976 -1 0 -270570
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_78
timestamp 1717613630
transform 0 1 34435 -1 0 -270573
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_79
timestamp 1717613630
transform 0 1 34426 -1 0 -271095
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_80
timestamp 1717613630
transform 0 1 33702 -1 0 -270969
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_81
timestamp 1717613630
transform 0 1 36791 -1 0 -270437
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_82
timestamp 1717613630
transform 0 1 36425 -1 0 -270433
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_83
timestamp 1717613630
transform 0 1 36256 -1 0 -270433
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_84
timestamp 1717613630
transform 0 1 35882 -1 0 -270433
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_85
timestamp 1717613630
transform 0 1 35713 -1 0 -270431
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_86
timestamp 1717613630
transform 0 1 35334 -1 0 -270428
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_87
timestamp 1717613630
transform 0 1 35164 -1 0 -270426
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_88
timestamp 1717613630
transform 0 1 34787 -1 0 -270413
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_89
timestamp 1717613630
transform 0 1 34619 -1 0 -270412
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_90
timestamp 1717613630
transform 0 1 34245 -1 0 -270400
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_91
timestamp 1717613630
transform 0 1 34610 -1 0 -270994
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_92
timestamp 1717613630
transform 0 1 34245 -1 0 -270975
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_93
timestamp 1717613630
transform 0 1 34077 -1 0 -270973
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_94
timestamp 1717613630
transform 0 1 37515 -1 0 -272141
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_95
timestamp 1717613630
transform 0 1 34324 -1 0 -271929
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_96
timestamp 1717613630
transform 0 1 36085 -1 0 -272142
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_97
timestamp 1717613630
transform 0 1 35647 -1 0 -272142
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_98
timestamp 1717613630
transform 0 1 36522 -1 0 -272141
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_99
timestamp 1717613630
transform 0 1 36296 -1 0 -271922
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_100
timestamp 1717613630
transform 0 1 35865 -1 0 -271925
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_101
timestamp 1717613630
transform 0 1 35427 -1 0 -271922
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_102
timestamp 1717613630
transform 0 1 35003 -1 0 -271922
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_103
timestamp 1717613630
transform 0 1 33890 -1 0 -271097
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_104
timestamp 1717613630
transform 0 1 31124 1 0 -300373
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_105
timestamp 1717613630
transform 0 1 32370 -1 0 -271375
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_106
timestamp 1717613630
transform 0 1 34586 -1 0 -271910
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_107
timestamp 1717613630
transform 0 1 31308 -1 0 -270785
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_108
timestamp 1717613630
transform 0 1 32840 -1 0 -270577
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_109
timestamp 1717613630
transform 0 1 32403 -1 0 -270580
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_110
timestamp 1717613630
transform 0 1 31966 -1 0 -270577
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_111
timestamp 1717613630
transform 0 1 31524 -1 0 -270580
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_112
timestamp 1717613630
transform 0 1 31090 -1 0 -270580
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_113
timestamp 1717613630
transform 0 1 31745 -1 0 -270791
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_114
timestamp 1717613630
transform 0 1 32611 -1 0 -270783
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_115
timestamp 1717613630
transform 0 1 32180 -1 0 -270787
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_116
timestamp 1717613630
transform 0 1 33198 1 0 -301396
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_117
timestamp 1717613630
transform 0 1 33201 1 0 -301026
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_118
timestamp 1717613630
transform 0 1 33212 1 0 -300373
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_119
timestamp 1717613630
transform 0 1 33105 1 0 -300370
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_120
timestamp 1717613630
transform 0 1 32997 1 0 -300372
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_121
timestamp 1717613630
transform 0 1 32789 1 0 -300372
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_122
timestamp 1717613630
transform 0 1 32686 1 0 -300372
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_123
timestamp 1717613630
transform 0 1 32478 1 0 -300372
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_124
timestamp 1717613630
transform -1 0 40130 0 1 -276637
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_125
timestamp 1717613630
transform 0 1 32164 1 0 -300372
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_126
timestamp 1717613630
transform 0 1 32039 1 0 -300373
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_127
timestamp 1717613630
transform 0 1 31852 1 0 -300361
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_128
timestamp 1717613630
transform 0 1 31713 1 0 -300368
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_129
timestamp 1717613630
transform 0 1 31600 1 0 -300368
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_130
timestamp 1717613630
transform 0 1 31367 1 0 -300368
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_131
timestamp 1717613630
transform 0 1 31251 1 0 -300370
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_132
timestamp 1717613630
transform 0 1 32969 1 0 -301024
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_133
timestamp 1717613630
transform 0 1 33086 1 0 -301387
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_134
timestamp 1717613630
transform 0 1 32976 1 0 -301387
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_135
timestamp 1717613630
transform 0 1 32141 1 0 -301385
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_136
timestamp 1717613630
transform 0 1 33084 1 0 -301022
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_137
timestamp 1717613630
transform 0 1 32782 1 0 -301016
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_138
timestamp 1717613630
transform 0 1 32660 1 0 -301016
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_139
timestamp 1717613630
transform 0 1 32650 1 0 -301394
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_140
timestamp 1717613630
transform 0 1 32780 1 0 -301394
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_141
timestamp 1717613630
transform 0 1 32468 1 0 -301392
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_142
timestamp 1717613630
transform 0 1 32336 1 0 -301390
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_143
timestamp 1717613630
transform 0 1 32341 1 0 -301021
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_144
timestamp 1717613630
transform 0 1 32468 1 0 -301021
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_145
timestamp 1717613630
transform 0 1 32155 1 0 -301021
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_146
timestamp 1717613630
transform 0 1 32025 1 0 -301017
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_147
timestamp 1717613630
transform 0 1 31229 1 0 -301054
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_148
timestamp 1717613630
transform 0 1 32018 1 0 -301387
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_149
timestamp 1717613630
transform 0 1 31730 1 0 -301484
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_150
timestamp 1717613630
transform 0 1 31565 1 0 -301486
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_151
timestamp 1717613630
transform 0 1 31378 1 0 -301486
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_152
timestamp 1717613630
transform 0 1 31220 1 0 -301484
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_153
timestamp 1717613630
transform 0 1 31716 1 0 -301050
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_154
timestamp 1717613630
transform 0 1 31376 1 0 -301052
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_155
timestamp 1717613630
transform 0 1 31581 1 0 -301048
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_156
timestamp 1717613630
transform 0 1 32358 1 0 -300373
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_157
timestamp 1717613630
transform -1 0 41095 0 1 -276631
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_158
timestamp 1717613630
transform -1 0 40793 0 1 -276629
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_159
timestamp 1717613630
transform -1 0 40485 0 1 -276631
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_160
timestamp 1717613630
transform 1 0 12480 0 1 -276586
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_161
timestamp 1717613630
transform 1 0 10958 0 1 -276553
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_162
timestamp 1717613630
transform 1 0 11684 0 1 -276750
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_163
timestamp 1717613630
transform 1 0 11758 0 1 -276649
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_164
timestamp 1717613630
transform 1 0 11211 0 1 -277277
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_165
timestamp 1717613630
transform 1 0 11484 0 1 -277849
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_166
timestamp 1717613630
transform 1 0 11929 0 1 -277275
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_167
timestamp 1717613630
transform 1 0 12192 0 1 -276638
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_168
timestamp 1717613630
transform 1 0 12186 0 1 -276835
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_169
timestamp 1717613630
transform 0 1 37685 -1 0 -268971
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_170
timestamp 1717613630
transform 0 1 37685 -1 0 -268424
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_171
timestamp 1717613630
transform 1 0 12471 0 1 -277355
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_172
timestamp 1717613630
transform 1 0 12192 0 1 -277261
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_173
timestamp 1717613630
transform 1 0 13609 0 1 -277692
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_174
timestamp 1717613630
transform 1 0 13492 0 1 -277925
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_175
timestamp 1717613630
transform 1 0 12193 0 1 -277923
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_176
timestamp 1717613630
transform 1 0 11697 0 1 -277772
box 16088 -7932 16222 -7868
use por_via_2cut  por_via_2cut_177
timestamp 1717613630
transform 0 1 38199 -1 0 -271021
box 16088 -7932 16222 -7868
use por_via_4cut  por_via_4cut_0
timestamp 1717613630
transform 1 0 15491 0 1 -279659
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_1
timestamp 1717613630
transform 1 0 16251 0 1 -279654
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_2
timestamp 1717613630
transform 1 0 15906 0 1 -279654
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_3
timestamp 1717613630
transform 1 0 14232 0 1 -279037
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_4
timestamp 1717613630
transform 0 1 37061 -1 0 -272147
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_5
timestamp 1717613630
transform 1 0 14260 0 1 -279828
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_6
timestamp 1717613630
transform 0 1 36877 -1 0 -270786
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_7
timestamp 1717613630
transform 0 1 36762 -1 0 -272168
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_8
timestamp 1717613630
transform -1 0 43094 0 -1 -295740
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_9
timestamp 1717613630
transform -1 0 44841 0 -1 -295507
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_10
timestamp 1717613630
transform -1 0 39210 0 -1 -295122
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_11
timestamp 1717613630
transform 0 1 31868 -1 0 -271608
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_12
timestamp 1717613630
transform 0 1 31641 -1 0 -271614
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_13
timestamp 1717613630
transform 0 1 31372 -1 0 -271556
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_14
timestamp 1717613630
transform 1 0 14257 0 1 -279646
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_15
timestamp 1717613630
transform 1 0 9448 0 1 -276623
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_16
timestamp 1717613630
transform 1 0 16689 0 1 -279648
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_17
timestamp 1717613630
transform 1 0 14671 0 1 -278888
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_18
timestamp 1717613630
transform -1 0 33617 0 -1 -294053
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_19
timestamp 1717613630
transform 1 0 14945 0 1 -279669
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_20
timestamp 1717613630
transform 1 0 15981 0 1 -280319
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_21
timestamp 1717613630
transform -1 0 45427 0 -1 -293841
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_22
timestamp 1717613630
transform -1 0 45357 0 -1 -295496
box 15948 -7932 16222 -7868
use sky130_fd_pr__cap_mim_m3_1_EEU5EF  sky130_fd_pr__cap_mim_m3_1_EEU5EF_0 paramcells
timestamp 1717613630
transform 0 -1 20303 -1 0 -279723
box -4192 -17600 3692 18302
use sky130_fd_pr__cap_mim_m3_1_EEU5EF  sky130_fd_pr__cap_mim_m3_1_EEU5EF_1
timestamp 1717613630
transform 0 -1 20294 1 0 -292633
box -4192 -17600 3692 18302
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_0 paramcells
timestamp 1717527227
transform -1 0 23102 0 1 -287324
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_1
timestamp 1717527227
transform -1 0 26798 0 1 -284831
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_2
timestamp 1717527227
transform -1 0 26755 0 1 -287330
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_RRZ644  sky130_fd_pr__cap_mim_m3_1_RRZ644_0 paramcells
timestamp 1717527227
transform -1 0 23271 0 1 -284613
box -986 -840 986 840
use sky130_fd_pr__cap_mim_m3_1_TBT74C  sky130_fd_pr__cap_mim_m3_1_TBT74C_0 paramcells
timestamp 1717527227
transform -1 0 36191 0 1 -286071
box -1786 -1640 1786 1640
use sky130_fd_pr__cap_mim_m3_1_TBT74C  sky130_fd_pr__cap_mim_m3_1_TBT74C_1
timestamp 1717527227
transform -1 0 19431 0 1 -286149
box -1786 -1640 1786 1640
use sky130_fd_pr__cap_mim_m3_1_TBT74C  sky130_fd_pr__cap_mim_m3_1_TBT74C_2
timestamp 1717527227
transform -1 0 31222 0 1 -286102
box -1786 -1640 1786 1640
use sky130_fd_pr__cap_mim_m3_2_2V27AY  sky130_fd_pr__cap_mim_m3_2_2V27AY_0 paramcells
timestamp 1717613630
transform 0 -1 19952 -1 0 -293305
box -4098 -18000 4120 18000
use sky130_fd_pr__cap_mim_m3_2_2V27AY  sky130_fd_pr__cap_mim_m3_2_2V27AY_1
timestamp 1717613630
transform 0 -1 19961 1 0 -279065
box -4098 -18000 4120 18000
use sky130_fd_pr__cap_mim_m3_2_4PHTN9  sky130_fd_pr__cap_mim_m3_2_4PHTN9_0 paramcells
timestamp 1717527227
transform 1 0 27164 0 1 -287318
box -1349 -1081 1371 1081
use sky130_fd_pr__cap_mim_m3_2_RQPX7Z  sky130_fd_pr__cap_mim_m3_2_RQPX7Z_0 paramcells
timestamp 1717527227
transform 1 0 36641 0 -1 -286081
box -1949 -1681 1971 1681
use sky130_fd_pr__pfet_01v8_XPC8Y6  sky130_fd_pr__pfet_01v8_XPC8Y6_1 paramcells
array 0 6 544 0 0 638
timestamp 1717527227
transform 1 0 26531 0 1 -286687
box -325 -319 325 319
use sky130_fd_pr__res_xhigh_po_0p69_KA8C77  sky130_fd_pr__res_xhigh_po_0p69_KA8C77_2 paramcells
timestamp 1717527227
transform 1 0 19503 0 1 -287933
box -2926 -1582 2926 1582
use sky130_fd_pr__res_xhigh_po_0p69_KA8C77  sky130_fd_pr__res_xhigh_po_0p69_KA8C77_3
timestamp 1717527227
transform 1 0 19502 0 1 -284399
box -2926 -1582 2926 1582
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 27235 0 1 -285414
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 27235 0 -1 -284326
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 27603 0 -1 -284326
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1715205430
transform 1 0 30179 0 1 -285414
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1715205430
transform 1 0 30179 0 -1 -284326
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 27695 0 -1 -284326
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 28339 0 1 -285414
box -38 -48 1878 592
use levelShifter  x3
timestamp 1717613630
transform 1 0 30687 0 1 -283596
box 609 -1772 4022 507
use TieH_1p8  x4
timestamp 1717613630
transform 1 0 25901 0 1 -284626
box 346 -837 1050 296
use sky130_fd_sc_hd__dfrtn_1  x5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 28339 0 -1 -284326
box -38 -48 1878 592
use sky130_fd_pr__cap_mim_m3_2_RQPX7Z  XC1
timestamp 1717527227
transform 1 0 19865 0 1 -286108
box -1949 -1681 1971 1681
use sky130_fd_pr__cap_mim_m3_2_HYMU45  XC3 paramcells
timestamp 1717527227
transform 1 0 23682 0 1 -284596
box -1149 -881 1171 881
use sky130_fd_pr__cap_mim_m3_2_4PHTN9  XC4
timestamp 1717527227
transform 1 0 23491 0 1 -287326
box -1349 -1081 1371 1081
use sky130_fd_pr__cap_mim_m3_2_RQPX7Z  XC5
timestamp 1717527227
transform 1 0 31657 0 -1 -286108
box -1949 -1681 1971 1681
use sky130_fd_pr__cap_mim_m3_2_4PHTN9  XC9
timestamp 1717527227
transform 1 0 27204 0 1 -284827
box -1349 -1081 1371 1081
use sky130_fd_pr__pfet_01v8_XPC8Y6  XM1
timestamp 1717527227
transform 1 0 25987 0 1 -287219
box -325 -319 325 319
use sky130_fd_pr__pfet_01v8_SKYQWJ  XM2 paramcells
timestamp 1717527227
transform 1 0 23405 0 -1 -285110
box -226 -537 226 537
use sky130_fd_pr__pfet_01v8_SKYQWJ  XM3
timestamp 1717527227
transform 1 0 23751 0 -1 -285110
box -226 -537 226 537
use sky130_fd_pr__nfet_01v8_5QNSAB  XM4 paramcells
timestamp 1717527227
transform 1 0 32643 0 1 -287844
box -263 -260 263 260
use sky130_fd_pr__nfet_01v8_G7LLWL  XM5 paramcells
timestamp 1717527227
transform 1 0 31469 0 1 -288426
box -285 -260 285 260
use sky130_fd_pr__nfet_01v8_G7LLWL  XM6
timestamp 1717527227
transform 1 0 31933 0 1 -288426
box -285 -260 285 260
use sky130_fd_pr__nfet_01v8_G7LLWL  XM7
timestamp 1717527227
transform 1 0 23352 0 -1 -284215
box -285 -260 285 260
use sky130_fd_pr__nfet_01v8_G7LLWL  XM8
timestamp 1717527227
transform 1 0 23816 0 -1 -284215
box -285 -260 285 260
use sky130_fd_pr__pfet_01v8_X6XW7S  XM9 paramcells
timestamp 1717527227
transform 1 0 32649 0 1 -287059
box -263 -477 263 477
use sky130_fd_pr__pfet_01v8_6QC8WZ  XM10 paramcells
timestamp 1717527227
transform 1 0 30399 0 1 -287219
box -285 -319 285 319
use sky130_fd_pr__pfet_g5v0d10v5_PQJ659  XM11 paramcells
timestamp 1717527227
transform 1 0 24088 0 1 -287669
box -338 -497 338 497
use sky130_fd_pr__pfet_01v8_GHZ9W9  XM12 paramcells
timestamp 1717527227
transform 1 0 30299 0 1 -286687
box -285 -319 285 319
use sky130_fd_pr__nfet_01v8_G7LLWL  XM13
timestamp 1717527227
transform 1 0 31465 0 1 -287844
box -285 -260 285 260
use sky130_fd_pr__pfet_01v8_SKYQWJ  XM14
timestamp 1717527227
transform 1 0 31170 0 1 -287001
box -226 -537 226 537
use sky130_fd_pr__pfet_01v8_XPC8Y6  XM16
timestamp 1717527227
transform 1 0 27075 0 1 -287219
box -325 -319 325 319
use sky130_fd_pr__nfet_g5v0d10v5_ESEQJ8  XM17 paramcells
timestamp 1717527227
transform 1 0 29004 0 1 -288194
box -318 -458 318 458
use sky130_fd_pr__pfet_g5v0d10v5_PQJ659  XM18
timestamp 1717527227
transform 1 0 24574 0 1 -287669
box -338 -497 338 497
use sky130_fd_pr__nfet_g5v0d10v5_SYBQJL  XM19 paramcells
timestamp 1717527227
transform 1 0 27854 0 1 -288194
box -962 -458 962 458
use sky130_fd_pr__pfet_01v8_XPC8Y6  XM20
timestamp 1717527227
transform 1 0 26531 0 1 -287219
box -325 -319 325 319
use sky130_fd_pr__nfet_g5v0d10v5_XSEQJ6  XM21 paramcells
timestamp 1717527227
transform 1 0 29827 0 1 -288194
box -635 -458 635 458
use sky130_fd_pr__pfet_01v8_XPC8Y6  XM22
array 0 3 544 0 0 640
timestamp 1717527227
transform 1 0 27619 0 1 -287219
box -325 -319 325 319
use sky130_fd_pr__pfet_01v8_XPC8Y6  XM23
timestamp 1717527227
transform 1 0 29795 0 1 -287219
box -325 -319 325 319
use sky130_fd_pr__pfet_g5v0d10v5_PQJ659  XM24
timestamp 1717527227
transform 1 0 23602 0 1 -287669
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_KLZS5A  XM25 paramcells
timestamp 1717527227
transform 1 0 24065 0 1 -286865
box -1101 -497 1101 497
use sky130_fd_pr__nfet_g5v0d10v5_69TNYL  XM26 paramcells
timestamp 1717527227
transform 1 0 26554 0 1 -288092
box -328 -358 328 358
use sky130_fd_pr__nfet_01v8_L9ESAD  XM27 paramcells
timestamp 1717527227
transform 1 0 31855 0 1 -287844
box -211 -260 211 260
use sky130_fd_pr__pfet_01v8_U6B66J  XM29 paramcells
timestamp 1717527227
transform 1 0 31861 0 1 -287059
box -211 -477 211 477
use sky130_fd_pr__nfet_01v8_5QNSAB  XM30
timestamp 1717527227
transform 1 0 32223 0 1 -287844
box -263 -260 263 260
use sky130_fd_pr__pfet_01v8_X6XW7S  XM31
timestamp 1717527227
transform 1 0 32229 0 1 -287059
box -263 -477 263 477
use sky130_fd_pr__nfet_01v8_L9ESAD  XM32
timestamp 1717527227
transform 1 0 24206 0 -1 -284215
box -211 -260 211 260
use sky130_fd_pr__pfet_01v8_U6B66J  XM33
timestamp 1717527227
transform 1 0 24188 0 -1 -285050
box -211 -477 211 477
use sky130_fd_pr__nfet_01v8_L9ESAD  XM34
timestamp 1717527227
transform 1 0 24522 0 -1 -284215
box -211 -260 211 260
use sky130_fd_pr__pfet_01v8_U6B66J  XM35
timestamp 1717527227
transform 1 0 24504 0 -1 -285050
box -211 -477 211 477
use sky130_fd_pr__nfet_01v8_5QNSAB  XM36
timestamp 1717527227
transform 1 0 25206 0 -1 -284215
box -263 -260 263 260
use sky130_fd_pr__nfet_01v8_L9ESAD  XM38
timestamp 1717527227
transform 1 0 24838 0 -1 -284215
box -211 -260 211 260
use sky130_fd_pr__pfet_01v8_U6B66J  XM39
timestamp 1717527227
transform 1 0 24820 0 -1 -285050
box -211 -477 211 477
use sky130_fd_pr__pfet_01v8_X6XW7S  XM40
timestamp 1717527227
transform 1 0 25188 0 -1 -285050
box -263 -477 263 477
<< labels >>
flabel metal1 27598 -287603 27598 -287603 0 FreeSans 400 0 0 0 vbp1
flabel metal1 29797 -287599 29797 -287599 0 FreeSans 400 0 0 0 vbp2
flabel metal1 29798 -287846 29798 -287846 0 FreeSans 400 0 0 0 vbn1
flabel metal1 30270 -287649 30270 -287649 0 FreeSans 400 0 0 0 VT2
flabel metal1 26133 -287918 26133 -287918 0 FreeSans 400 0 0 0 Vbg
flabel metal1 31004 -287558 31004 -287558 0 FreeSans 400 0 0 0 VT3
flabel metal2 32747 -287555 32747 -287555 0 FreeSans 400 0 0 0 Td_Lb
flabel metal2 32334 -287557 32334 -287557 0 FreeSans 400 0 0 0 Td_L
flabel metal2 32599 -288423 32599 -288423 0 FreeSans 400 0 0 0 VSS
flabel metal2 32417 -286352 32417 -286352 0 FreeSans 400 0 0 0 VCCL
flabel metal2 25218 -286723 25218 -286723 0 FreeSans 400 0 0 0 VCCH
flabel metal1 23057 -284645 23057 -284645 0 FreeSans 400 0 0 0 din
flabel metal2 23807 -284534 23807 -284534 0 FreeSans 400 0 0 0 Td_S
flabel metal2 25245 -284524 25245 -284524 0 FreeSans 400 0 0 0 Td_Sd
flabel metal2 24391 -285633 24391 -285633 0 FreeSans 400 0 0 0 VCCL
flabel metal2 24417 -283903 24417 -283903 0 FreeSans 400 0 0 0 VSS
flabel metal2 36799 -284322 36799 -284322 0 FreeSans 400 0 0 0 porb_h
flabel metal2 16520 -286264 16720 -286064 0 FreeSans 256 0 0 0 din
port 0 nsew
flabel metal2 36783 -286341 36783 -286341 0 FreeSans 400 0 0 0 porb
flabel metal2 30469 -283777 30669 -283577 0 FreeSans 256 0 0 0 VCCL
port 2 nsew
flabel metal2 36711 -288173 36815 -288112 0 FreeSans 400 0 0 0 por
flabel metal2 36844 -284387 37044 -284187 0 FreeSans 256 0 0 0 porb_h
port 7 nsew
flabel metal2 36830 -286437 37030 -286237 0 FreeSans 256 0 0 0 porb
port 6 nsew
flabel metal2 36815 -288245 37015 -288045 0 FreeSans 256 0 0 0 por
port 1 nsew
flabel metal1 30961 -284690 30961 -284690 0 FreeSans 400 0 0 0 porbPre
flabel metal1 30961 -285019 30961 -285019 0 FreeSans 400 0 0 0 porPre
flabel metal2 23866 -288669 24066 -288469 0 FreeSans 256 0 0 0 VSS
port 3 nsew
flabel metal1 16345 -289669 16545 -289469 0 FreeSans 256 0 0 0 Vbg
port 4 nsew
<< end >>
