magic
tech sky130A
magscale 1 2
timestamp 1717527227
<< pwell >>
rect -515 -358 515 358
<< mvnmos >>
rect -287 -100 -187 100
rect -129 -100 -29 100
rect 29 -100 129 100
rect 187 -100 287 100
<< mvndiff >>
rect -345 88 -287 100
rect -345 -88 -333 88
rect -299 -88 -287 88
rect -345 -100 -287 -88
rect -187 88 -129 100
rect -187 -88 -175 88
rect -141 -88 -129 88
rect -187 -100 -129 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 129 88 187 100
rect 129 -88 141 88
rect 175 -88 187 88
rect 129 -100 187 -88
rect 287 88 345 100
rect 287 -88 299 88
rect 333 -88 345 88
rect 287 -100 345 -88
<< mvndiffc >>
rect -333 -88 -299 88
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect 299 -88 333 88
<< mvpsubdiff >>
rect -479 310 479 322
rect -479 276 -371 310
rect 371 276 479 310
rect -479 264 479 276
rect -479 214 -421 264
rect -479 -214 -467 214
rect -433 -214 -421 214
rect 421 214 479 264
rect -479 -264 -421 -214
rect 421 -214 433 214
rect 467 -214 479 214
rect 421 -264 479 -214
rect -479 -276 479 -264
rect -479 -310 -371 -276
rect 371 -310 479 -276
rect -479 -322 479 -310
<< mvpsubdiffcont >>
rect -371 276 371 310
rect -467 -214 -433 214
rect 433 -214 467 214
rect -371 -310 371 -276
<< poly >>
rect -287 172 -187 188
rect -287 138 -271 172
rect -203 138 -187 172
rect -287 100 -187 138
rect -129 172 -29 188
rect -129 138 -113 172
rect -45 138 -29 172
rect -129 100 -29 138
rect 29 172 129 188
rect 29 138 45 172
rect 113 138 129 172
rect 29 100 129 138
rect 187 172 287 188
rect 187 138 203 172
rect 271 138 287 172
rect 187 100 287 138
rect -287 -138 -187 -100
rect -287 -172 -271 -138
rect -203 -172 -187 -138
rect -287 -188 -187 -172
rect -129 -138 -29 -100
rect -129 -172 -113 -138
rect -45 -172 -29 -138
rect -129 -188 -29 -172
rect 29 -138 129 -100
rect 29 -172 45 -138
rect 113 -172 129 -138
rect 29 -188 129 -172
rect 187 -138 287 -100
rect 187 -172 203 -138
rect 271 -172 287 -138
rect 187 -188 287 -172
<< polycont >>
rect -271 138 -203 172
rect -113 138 -45 172
rect 45 138 113 172
rect 203 138 271 172
rect -271 -172 -203 -138
rect -113 -172 -45 -138
rect 45 -172 113 -138
rect 203 -172 271 -138
<< locali >>
rect -467 276 -371 310
rect 371 276 467 310
rect -467 214 -433 276
rect 433 214 467 276
rect -287 138 -271 172
rect -203 138 -187 172
rect -129 138 -113 172
rect -45 138 -29 172
rect 29 138 45 172
rect 113 138 129 172
rect 187 138 203 172
rect 271 138 287 172
rect -333 88 -299 104
rect -333 -104 -299 -88
rect -175 88 -141 104
rect -175 -104 -141 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 141 88 175 104
rect 141 -104 175 -88
rect 299 88 333 104
rect 299 -104 333 -88
rect -287 -172 -271 -138
rect -203 -172 -187 -138
rect -129 -172 -113 -138
rect -45 -172 -29 -138
rect 29 -172 45 -138
rect 113 -172 129 -138
rect 187 -172 203 -138
rect 271 -172 287 -138
rect -467 -276 -433 -214
rect 433 -276 467 -214
rect -467 -310 -371 -276
rect 371 -310 467 -276
<< viali >>
rect -271 138 -203 172
rect -113 138 -45 172
rect 45 138 113 172
rect 203 138 271 172
rect -333 -88 -299 88
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect 299 -88 333 88
rect -271 -172 -203 -138
rect -113 -172 -45 -138
rect 45 -172 113 -138
rect 203 -172 271 -138
<< metal1 >>
rect -283 172 -191 178
rect -283 138 -271 172
rect -203 138 -191 172
rect -283 132 -191 138
rect -125 172 -33 178
rect -125 138 -113 172
rect -45 138 -33 172
rect -125 132 -33 138
rect 33 172 125 178
rect 33 138 45 172
rect 113 138 125 172
rect 33 132 125 138
rect 191 172 283 178
rect 191 138 203 172
rect 271 138 283 172
rect 191 132 283 138
rect -339 88 -293 100
rect -339 -88 -333 88
rect -299 -88 -293 88
rect -339 -100 -293 -88
rect -181 88 -135 100
rect -181 -88 -175 88
rect -141 -88 -135 88
rect -181 -100 -135 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 135 88 181 100
rect 135 -88 141 88
rect 175 -88 181 88
rect 135 -100 181 -88
rect 293 88 339 100
rect 293 -88 299 88
rect 333 -88 339 88
rect 293 -100 339 -88
rect -283 -138 -191 -132
rect -283 -172 -271 -138
rect -203 -172 -191 -138
rect -283 -178 -191 -172
rect -125 -138 -33 -132
rect -125 -172 -113 -138
rect -45 -172 -33 -138
rect -125 -178 -33 -172
rect 33 -138 125 -132
rect 33 -172 45 -138
rect 113 -172 125 -138
rect 33 -178 125 -172
rect 191 -138 283 -132
rect 191 -172 203 -138
rect 271 -172 283 -138
rect 191 -178 283 -172
<< properties >>
string FIXED_BBOX -450 -293 450 293
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1 l 0.50 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
