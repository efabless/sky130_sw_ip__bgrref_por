* NGSPICE file created from sky130_sw_ip__bgrref_por.ext - technology: sky130A

.subckt sky130_sw_ip__bgrref_por vbg por avss avdd dvdd porb dvss porb_h[0] porb_h[1]
X0 dvss.t440 x2.VT2.t0 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X1 dvss.t441 x2.VT3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X2 a_35262_n291454.t5 a_35074_n291454# dvdd.t285 dvdd.t283 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X3 a_29895_n287373# x2.Td_Sd.t6 dvdd.t170 dvdd.t169 sky130_fd_pr__pfet_01v8_hvt ad=0.1218 pd=1.42 as=0.07245 ps=0.765 w=0.42 l=0.15
X4 x2.Td_Sd.t0 a_25883_n288267.t4 dvdd.t274 dvdd.t273 sky130_fd_pr__pfet_01v8 ad=0.217 pd=2.02 as=0.1155 ps=1.03 w=0.7 l=0.15
X5 dvdd.t172 x2.Td_Sd.t7 a_29214_n287320# dvdd.t171 sky130_fd_pr__pfet_01v8_hvt ad=0.172775 pd=1.58 as=0.063 ps=0.72 w=0.42 l=0.15
X6 a_37002_n287783.t1 a_36398_n287783.t4 dvss.t108 dvss.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X7 x2.Td_L.t5 a_32918_n290853.t3 dvdd.t72 dvdd.t17 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.217 ps=2.02 w=0.7 l=0.15
X8 a_5972_n290308.t2 a_4566_n291516.t3 x1.vbn.t3 avss.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
X9 avdd.t77 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t4 porb_h[0].t22 avdd.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X10 a_25567_n288267.t3 a_25251_n288267.t4 dvdd.t181 dvdd.t180 sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.98 as=0.203 ps=1.98 w=0.7 l=0.15
X11 porb_h[1].t15 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t5 dvss.t71 dvss.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X12 a_29211_n288416# x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtp_1_0.D dvdd.t328 dvdd.t327 sky130_fd_pr__pfet_01v8_hvt ad=0.05985 pd=0.705 as=0.1197 ps=1.41 w=0.42 l=0.15
X13 avdd.t120 a_34073_n287091.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X14 a_30814_n289746# x2.vbp2 a_30112_n289746# dvdd.t12 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X15 a_32918_n290853.t0 a_32248_n290278# dvss.t204 dvss.t203 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
X16 a_18961_n289908# a_19195_n292308# dvss.t315 sky130_fd_pr__res_xhigh_po_0p69 l=10
X17 dvss.t261 x2.Td_Lb a_30075_n288356# dvss.t260 sky130_fd_pr__nfet_01v8 ad=0.211225 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X18 por.t47 a_35454_n291454.t24 dvdd.t81 dvdd.t51 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X19 dvdd.t119 x2.vbp1.t31 a_30112_n289746# dvdd.t11 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X20 a_30837_n288413# x2.Td_Lb dvss.t259 dvss.t258 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X21 por.t46 a_35454_n291454.t25 dvdd.t83 dvdd.t82 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X22 a_8490_n290308# a_8656_n292108# avss.t25 sky130_fd_pr__res_xhigh_po_0p35 l=7
X23 porb_h[0].t15 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t6 dvss.t318 dvss.t317 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X24 a_19662_n286374# a_19896_n288774# dvss.t177 sky130_fd_pr__res_xhigh_po_0p69 l=10
X25 a_29895_n287373# a_29481_n287384# a_29214_n287320# dvdd.t111 sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X26 a_29966_n288037# a_29487_n288398# a_29876_n288037# dvdd.t214 sky130_fd_pr__pfet_01v8_hvt ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X27 x2.VT3 x2.VT2.t8 a_30410_n291353# dvss.t125 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.3
X28 dvdd.t143 x2.vbp1.t32 a_28094_n290278.t7 dvdd.t43 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X29 a_34073_n287091.t3 x2.x3.S1B dvss.t13 dvss.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=0.5
X30 dvss.t442 x2.VT2.t3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X31 avdd.t95 x1.vt.t3 x1.vo.t2 avdd.t94 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
X32 porb.t15 a_35469_n289052.t24 dvss.t169 dvss.t168 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X33 dvss.t443 x2.VT2.t2 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X34 dvss.t366 x2.VT3 a_32248_n290278# dvss.t365 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.3
X35 a_9100_n286429# a_9266_n288829# avss.t55 sky130_fd_pr__res_xhigh_po_0p35 l=10
X36 dvss.t444 x2.VT2.t3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X37 a_35277_n289052.t5 a_35089_n289052# dvdd.t191 dvdd.t188 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X38 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtp_1_0.D a_27214_n288191# dvdd.t210 dvdd.t209 sky130_fd_pr__pfet_01v8 ad=0.0825 pd=0.83 as=0.155 ps=1.62 w=0.5 l=0.15
X39 dvss.t445 x2.VT2.t0 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X40 a_35469_n289052.t20 a_35277_n289052.t6 dvdd.t340 dvdd.t205 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X41 a_19662_n286374# a_19428_n288774# dvss.t85 sky130_fd_pr__res_xhigh_po_0p69 l=10
X42 dvss.t156 a_28056_n288420# x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N dvss.t155 sky130_fd_pr__nfet_01v8 ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X43 por.t15 a_35454_n291454.t26 dvss.t302 dvss.t301 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X44 dvdd.t239 a_35262_n291454.t6 a_35454_n291454.t23 dvdd.t231 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X45 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N a_28056_n288420# dvss.t154 dvss.t153 sky130_fd_pr__nfet_01v8 ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X46 x2.VT3 dvss.t364 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X47 x2.VT2.t0 dvss.t198 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X48 porb.t47 a_35469_n289052.t25 dvdd.t163 dvdd.t162 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X49 dvdd.t256 a_35454_n291454.t27 por.t45 dvdd.t255 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X50 dvss.t215 a_35089_n289052# a_35277_n289052.t1 dvss.t214 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X51 dvdd.t167 a_35469_n289052.t26 porb.t46 dvdd.t73 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X52 a_28094_n290278.t9 x2.vbp2 w_31992_n290497# dvdd.t14 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X53 dvdd.t235 a_35262_n291454.t7 a_35454_n291454.t22 dvdd.t92 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X54 dvss.t446 x2.VT3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X55 dvss.t76 a_37002_n287783.t4 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t1 dvss.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X56 a_8490_n290308# a_7996_n292010# avss.t0 sky130_fd_pr__res_xhigh_po_0p35 l=7
X57 dvss.t190 a_35469_n289052.t27 porb.t14 dvss.t189 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X58 x2.VT3 dvss.t363 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X59 x2.VT2.t3 dvss.t329 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X60 a_9764_n286429# a_9930_n288829# avss.t54 sky130_fd_pr__res_xhigh_po_0p35 l=10
X61 a_25567_n288267.t0 dvss.t207 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X62 dvdd.t139 a_35454_n291454.t28 por.t44 dvdd.t138 sky130_fd_pr__pfet_01v8 ad=0.217 pd=2.02 as=0.1155 ps=1.03 w=0.7 l=0.15
X63 a_11424_n286429# x1.Vinn.t0 avss.t31 sky130_fd_pr__res_xhigh_po_0p35 l=10
X64 a_18258_n286374# a_18024_n288774# dvss.t436 sky130_fd_pr__res_xhigh_po_0p69 l=10
X65 a_24270_n290121.t17 a_24270_n290121.t16 avdd.t5 avdd.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X66 a_8768_n286429# a_8934_n288829# avss.t24 sky130_fd_pr__res_xhigh_po_0p35 l=10
X67 dvdd.t341 a_35277_n289052.t7 a_35469_n289052.t21 dvdd.t311 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X68 porb_h[1].t31 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t7 avdd.t76 avdd.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X69 a_10428_n286429# a_10594_n288829# avss.t62 sky130_fd_pr__res_xhigh_po_0p35 l=10
X70 x2.VT2.t2 dvss.t333 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X71 porb_h[1].t30 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t8 avdd.t75 avdd.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X72 a_34073_n287091.t0 a_34015_n286994.t4 avdd.t1 avdd.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.841 pd=6.38 as=0.4205 ps=3.19 w=2.9 l=0.5
X73 dvdd.t324 a_15914_n289870# x2.din dvdd.t323 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X74 a_7772_n286429# a_7938_n288829# avss.t39 sky130_fd_pr__res_xhigh_po_0p35 l=10
X75 a_30410_n291353# x2.vbn1.t16 dvss.t423 dvss.t422 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.8
X76 dvss.t139 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t9 porb_h[1].t14 dvss.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X77 dvdd.t140 a_35454_n291454.t29 por.t43 dvdd.t84 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X78 dvss.t447 x2.VT3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X79 dvss.t382 a_35469_n289052.t28 porb.t13 dvss.t381 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X80 dvdd.t276 a_25883_n288267.t5 x2.Td_Sd.t1 dvdd.t275 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.217 ps=2.02 w=0.7 l=0.15
X81 dvdd.t62 x2.x3.S1 x2.x3.S1B dvdd.t61 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.217 ps=2.02 w=0.7 l=0.15
X82 a_30103_n287373# a_30022_n287538# a_30031_n287373# dvss.t236 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X83 avdd.t112 a_13449_n292106.t3 x1.vt.t2 avdd.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
X84 a_17790_n286374# a_18024_n288774# dvss.t435 sky130_fd_pr__res_xhigh_po_0p69 l=10
X85 a_17790_n286374# a_17790_n288774# dvss.t63 sky130_fd_pr__res_xhigh_po_0p69 l=10
X86 avdd.t79 x2.x3.aout.t3 a_36398_n287783.t0 avdd.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.58 as=0.3625 ps=2.79 w=2.5 l=0.5
X87 x2.VT2.t1 dvss.t418 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X88 dvdd.t193 a_35277_n289052.t8 a_35469_n289052.t8 dvdd.t192 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X89 x2.vbp1.t27 x2.vbp1.t26 dvdd.t155 dvdd.t154 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X90 dvss.t448 x2.VT3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X91 dvdd.t196 a_35454_n291454.t30 por.t42 dvdd.t195 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X92 a_13144_n286429# a_13310_n288829# avss.t68 sky130_fd_pr__res_xhigh_po_0p35 l=10
X93 avdd.t70 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t10 porb_h[1].t29 avdd.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X94 a_29481_n287384# x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N dvss.t167 dvss.t166 sky130_fd_pr__nfet_01v8 ad=0.2035 pd=2.03 as=0.1212 ps=1.1 w=0.74 l=0.15
X95 dvdd.t294 a_35469_n289052.t29 porb.t45 dvdd.t265 sky130_fd_pr__pfet_01v8 ad=0.217 pd=2.02 as=0.1155 ps=1.03 w=0.7 l=0.15
X96 a_22470_n286374# a_22236_n288774# dvss.t9 sky130_fd_pr__res_xhigh_po_0p69 l=10
X97 a_35469_n289052.t9 a_35277_n289052.t9 dvss.t221 dvss.t220 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X98 x1.VD.t5 x1.Vinn.t2 x1.VS avss.t19 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X99 a_35454_n291454.t7 a_35262_n291454.t8 dvss.t276 dvss.t275 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X100 x1.VD.t4 x1.Vinn.t3 x1.VS avss.t20 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X101 a_29997_n288356# a_29671_n288104# a_29876_n288037# dvss.t264 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X102 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N a_28056_n288420# dvdd.t137 dvdd.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X103 a_30649_n288001# a_29671_n288104# a_30447_n288420# dvdd.t223 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X104 dvss.t184 x2.vbn1.t13 x2.vbn1.t14 dvss.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.8
X105 a_7772_n286429# a_7606_n288829# avss.t58 sky130_fd_pr__res_xhigh_po_0p35 l=10
X106 por.t14 a_35454_n291454.t31 dvss.t231 dvss.t230 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X107 dvdd.t190 a_35089_n289052# a_35277_n289052.t4 dvdd.t186 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X108 porb_h[1].t28 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t11 avdd.t74 avdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X109 a_28607_n287397# x2.Td_Sd.t8 a_28571_n287754# dvdd.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X110 x2.delayPulse_digital_0/sky130_fd_sc_ls__xor2_1_0.X a_28607_n287397# a_28768_n287754# dvdd.t164 sky130_fd_pr__pfet_01v8_hvt ad=0.3864 pd=2.93 as=0.196 ps=1.47 w=1.12 l=0.15
X111 dvdd.t157 x2.vbp1.t24 x2.vbp1.t25 dvdd.t156 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X112 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N a_28056_n288420# dvss.t152 dvss.t151 sky130_fd_pr__nfet_01v8 ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X113 avss.t11 x1.vbn.t4 x1.vo.t1 avss.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X114 dvss.t176 a_28607_n287397# x2.delayPulse_digital_0/sky130_fd_sc_ls__xor2_1_0.X dvss.t175 sky130_fd_pr__nfet_01v8 ad=0.2997 pd=2.29 as=0.1554 ps=1.16 w=0.74 l=0.15
X115 dvdd.t30 a_35469_n289052.t30 porb.t44 dvdd.t29 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X116 x2.vbp1.t23 x2.vbp1.t22 dvdd.t34 dvdd.t33 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X117 porb_h[0].t14 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t12 dvss.t67 dvss.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X118 porb_h[0].t13 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t13 dvss.t69 dvss.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X119 dvdd.t32 a_35469_n289052.t31 porb.t43 dvdd.t31 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X120 a_21066_n286374# a_20832_n288774# dvss.t62 sky130_fd_pr__res_xhigh_po_0p69 l=10
X121 por.t41 a_35454_n291454.t32 dvdd.t258 dvdd.t257 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X122 x2.x3.aout.t2 a_34073_n287091.t5 avdd.t81 avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.841 pd=6.38 as=0.4205 ps=3.19 w=2.9 l=0.5
X123 a_25883_n288267.t1 a_25567_n288267.t4 dvdd.t4 dvdd.t3 sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.98 as=0.203 ps=1.98 w=0.7 l=0.15
X124 avdd.t121 a_24270_n290121.t0 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X125 dvss.t408 a_24253_n287224.t4 x2.VT2.t6 dvss.t407 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.3
X126 porb_h[0].t27 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t14 avdd.t73 avdd.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X127 porb.t12 a_35469_n289052.t32 dvss.t36 dvss.t35 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X128 dvss.t78 a_32918_n290853.t4 x2.Td_L.t1 dvss.t77 sky130_fd_pr__nfet_01v8 ad=0.155 pd=1.62 as=0.0825 ps=0.83 w=0.5 l=0.15
X129 x2.Td_Lb x2.Td_L.t6 dvdd.t346 dvdd.t106 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.217 ps=2.02 w=0.7 l=0.15
X130 x2.VT3 x2.VT2.t9 dvdd.t290 dvdd.t289 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X131 por.t13 a_35454_n291454.t33 dvss.t304 dvss.t303 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X132 por.t40 a_35454_n291454.t34 dvdd.t342 dvdd.t112 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X133 a_34015_n286994.t1 x2.x3.S1 dvss.t53 dvss.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=0.5
X134 x2.VT2.t7 a_24253_n287224.t5 a_30814_n289746# dvdd.t320 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X135 dvdd.t121 a_30779_n287655# a_30728_n287754# dvdd.t120 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X136 a_18493_n289908# a_18259_n292308# dvss.t409 sky130_fd_pr__res_xhigh_po_0p69 l=10
X137 a_35469_n289052.t2 a_35277_n289052.t10 dvdd.t26 dvdd.t25 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X138 a_19194_n286374# a_19428_n288774# dvss.t249 sky130_fd_pr__res_xhigh_po_0p69 l=10
X139 a_34015_n286994.t3 a_34073_n287091.t6 avdd.t89 avdd.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0.841 pd=6.38 as=0.4205 ps=3.19 w=2.9 l=0.5
X140 dvss.t449 x2.VT3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X141 x2.VT3 dvss.t362 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X142 dvss.t278 a_35262_n291454.t9 a_35454_n291454.t6 dvss.t277 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X143 a_25251_n288267.t1 x2.Td_S.t4 dvdd.t50 dvdd.t49 sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.98 as=0.203 ps=1.98 w=0.7 l=0.15
X144 dvss.t33 x2.Td_Sd.t9 a_30103_n287373# dvss.t32 sky130_fd_pr__nfet_01v8 ad=0.240325 pd=1.715 as=0.0441 ps=0.63 w=0.42 l=0.15
X145 porb.t42 a_35469_n289052.t33 dvdd.t39 dvdd.t38 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X146 dvdd.t279 x2.vbp1.t20 x2.vbp1.t21 dvdd.t184 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X147 avdd.t72 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t15 porb_h[0].t26 avdd.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X148 x2.vbn1.t12 x2.vbn1.t11 dvss.t229 dvss.t228 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X149 a_23173_n289908# a_22939_n292308# dvss.t248 sky130_fd_pr__res_xhigh_po_0p69 l=10
X150 avdd.t71 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t16 porb_h[0].t28 avdd.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X151 dvss.t450 x2.VT3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X152 a_29688_n287709# a_29481_n287384# dvss.t114 dvss.t113 sky130_fd_pr__nfet_01v8 ad=0.2479 pd=2.15 as=0.3299 ps=2.67 w=0.74 l=0.15
X153 a_35469_n289052.t3 a_35277_n289052.t11 dvdd.t28 dvdd.t27 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X154 a_18726_n286374# a_18960_n288774# dvss.t247 sky130_fd_pr__res_xhigh_po_0p69 l=10
X155 dvss.t122 a_36398_n287783.t5 a_37002_n287783.t0 dvss.t121 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X156 porb.t11 a_35469_n289052.t34 dvss.t41 dvss.t40 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X157 porb.t41 a_35469_n289052.t35 dvdd.t46 dvdd.t45 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X158 dvdd.t37 x2.Td_Sd.t10 a_29487_n288398# dvdd.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.31 ps=2.62 w=1 l=0.15
X159 a_14140_n286429# a_14306_n288829# avss.t30 sky130_fd_pr__res_xhigh_po_0p35 l=10
X160 x2.VT3 dvss.t361 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X161 avdd.t69 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t17 porb_h[1].t27 avdd.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X162 dvdd.t243 a_31045_n288085# x2.porPre dvdd.t242 sky130_fd_pr__pfet_01v8_hvt ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X163 x2.porbPre a_31115_n287366# dvss.t161 dvss.t160 sky130_fd_pr__nfet_01v8 ad=0.2146 pd=2.06 as=0.126075 ps=1.1 w=0.74 l=0.15
X164 dvdd.t44 x2.vbp1.t18 x2.vbp1.t19 dvdd.t43 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X165 dvss.t451 x2.VT2.t3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X166 a_25567_n288267.t2 a_25251_n288267.t5 dvdd.t182 dvdd.t180 sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.98 as=0.203 ps=1.98 w=0.7 l=0.15
X167 dvss.t434 a_35454_n291454.t35 por.t12 dvss.t433 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X168 a_35262_n291454.t4 a_35074_n291454# dvdd.t284 dvdd.t283 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X169 dvss.t65 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t18 porb_h[0].t12 dvss.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0.2025 pd=2.04 as=0.105 ps=1.03 w=0.75 l=0.5
X170 a_9764_n286429# a_9598_n288829# avss.t22 sky130_fd_pr__res_xhigh_po_0p35 l=10
X171 dvdd.t345 a_35277_n289052.t12 a_35469_n289052.t22 dvdd.t77 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X172 avss.t10 x1.vbn.t5 x1.vo.t0 avss.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X173 a_31045_n288085# a_30447_n288420# dvss.t292 dvss.t291 sky130_fd_pr__nfet_01v8 ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X174 a_8768_n286429# a_8602_n288829# avss.t57 sky130_fd_pr__res_xhigh_po_0p35 l=10
X175 dvss.t452 x2.VT2.t3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X176 por.t39 a_35454_n291454.t36 dvdd.t52 dvdd.t51 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X177 porb.t40 a_35469_n289052.t36 dvdd.t114 dvdd.t100 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X178 a_35454_n291454.t21 a_35262_n291454.t10 dvdd.t91 dvdd.t90 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X179 porb_h[1].t13 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t19 dvss.t294 dvss.t293 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X180 a_29998_n287709# a_29688_n287709# a_29895_n287373# dvdd.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X181 a_19897_n289908# a_19663_n292308# dvss.t279 sky130_fd_pr__res_xhigh_po_0p69 l=10
X182 a_22002_n286374# a_22236_n288774# dvss.t342 sky130_fd_pr__res_xhigh_po_0p69 l=10
X183 a_28571_n287754# x2.Td_L.t7 dvdd.t348 dvdd.t347 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X184 porb_h[0].t11 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t20 dvss.t296 dvss.t295 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X185 porb_h[0].t10 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t21 dvss.t223 dvss.t222 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X186 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N a_28056_n288420# dvdd.t135 dvdd.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.435 as=0.1876 ps=1.455 w=1.12 l=0.15
X187 a_30112_n289746# x2.vbp2 a_30814_n289746# dvdd.t14 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X188 por.t38 a_35454_n291454.t37 dvdd.t54 dvdd.t53 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X189 a_14140_n286429# a_13974_n288829# avss.t61 sky130_fd_pr__res_xhigh_po_0p35 l=10
X190 a_24570_n290925.t3 a_24570_n290925.t2 a_24270_n290121.t1 avdd.t96 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
X191 a_13144_n286429# a_12978_n288829# avss.t60 sky130_fd_pr__res_xhigh_po_0p35 l=10
X192 x2.VT3 dvss.t360 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X193 dvss.t15 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t22 porb_h[1].t12 dvss.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X194 a_29876_n288037# x2.Td_Lb dvdd.t220 dvdd.t219 sky130_fd_pr__pfet_01v8_hvt ad=0.1239 pd=1.43 as=0.137125 ps=1.155 w=0.42 l=0.15
X195 x2.VT2.t0 dvss.t197 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X196 dvss.t453 x2.VT2.t1 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X197 a_19429_n289908# a_19663_n292308# dvss.t339 sky130_fd_pr__res_xhigh_po_0p69 l=10
X198 x1.Vinp.t1 x1.Vinn.t1 avss.t59 sky130_fd_pr__res_xhigh_po_0p35 l=9
X199 a_24270_n290121.t15 a_24270_n290121.t14 avdd.t83 avdd.t82 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X200 a_22002_n286374# a_21768_n288774# dvss.t367 sky130_fd_pr__res_xhigh_po_0p69 l=10
X201 x2.vbn1.t0 dvss.t170 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X202 dvss.t17 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t23 porb_h[0].t9 dvss.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X203 avdd.t19 avdd.t18 a_14970_n288829# avss.t15 sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.9
X204 a_20598_n286374# a_20364_n288774# dvss.t338 sky130_fd_pr__res_xhigh_po_0p69 l=10
X205 dvss.t454 x2.VT2.t3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X206 porb.t39 a_35469_n289052.t37 dvdd.t115 dvdd.t57 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X207 por.t37 a_35454_n291454.t38 dvdd.t296 dvdd.t295 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X208 dvdd.t93 a_35262_n291454.t11 a_35454_n291454.t20 dvdd.t92 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X209 x2.VT2.t3 dvss.t328 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X210 x2.x3.S1 x2.porbPre dvdd.t309 dvdd.t308 sky130_fd_pr__pfet_01v8 ad=0.217 pd=2.02 as=0.1155 ps=1.03 w=0.7 l=0.15
X211 a_28094_n290278.t6 x2.vbp1.t33 dvdd.t145 dvdd.t144 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X212 a_4566_n290308.t0 a_4508_n291419.t0 a_4508_n291419.t1 avdd.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X213 dvss.t439 a_35277_n289052.t13 a_35469_n289052.t23 dvss.t438 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X214 dvdd.t297 a_35454_n291454.t39 por.t36 dvdd.t138 sky130_fd_pr__pfet_01v8 ad=0.217 pd=2.02 as=0.1155 ps=1.03 w=0.7 l=0.15
X215 dvss.t235 x2.porPre a_35074_n291454# dvss.t234 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.155 ps=1.62 w=0.5 l=0.15
X216 dvdd.t95 a_35262_n291454.t12 a_35454_n291454.t19 dvdd.t94 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X217 a_18025_n289908# a_18259_n292308# dvss.t173 sky130_fd_pr__res_xhigh_po_0p69 l=10
X218 dvss.t402 a_24253_n287224.t6 x2.Td_S.t1 dvss.t401 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.3
X219 a_20130_n286374# a_20364_n288774# dvss.t437 sky130_fd_pr__res_xhigh_po_0p69 l=10
X220 dvss.t455 x2.VT3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X221 a_12812_n286429# a_12646_n288829# avss.t27 sky130_fd_pr__res_xhigh_po_0p35 l=10
X222 porb_h[0].t8 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t24 dvss.t26 dvss.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X223 dvss.t43 a_35469_n289052.t38 porb.t10 dvss.t42 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X224 dvss.t233 a_35454_n291454.t40 por.t11 dvss.t232 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X225 dvdd.t277 a_25883_n288267.t6 x2.Td_Sd.t2 dvdd.t275 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.217 ps=2.02 w=0.7 l=0.15
X226 a_30917_n287365# x2.Td_Sd.t11 dvss.t82 dvss.t81 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.0819 ps=0.81 w=0.42 l=0.15
X227 dvss.t456 x2.VT3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X228 a_32248_n290278# x2.VT3 w_31992_n290497# w_31992_n290497# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X229 dvdd.t48 a_35469_n289052.t39 porb.t38 dvdd.t47 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X230 dvss.t225 x2.vbn1.t9 x2.vbn1.t10 dvss.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X231 a_30011_n288135# a_29876_n288037# dvss.t431 dvss.t430 sky130_fd_pr__nfet_01v8 ad=0.24605 pd=1.405 as=0.211225 ps=1.45 w=0.74 l=0.15
X232 a_18025_n289908# a_17791_n292308# dvss.t4 sky130_fd_pr__res_xhigh_po_0p69 l=10
X233 a_17790_n288774# a_17791_n292308# dvss.t117 sky130_fd_pr__res_xhigh_po_0p69 l=10
X234 a_20130_n286374# a_19896_n288774# dvss.t178 sky130_fd_pr__res_xhigh_po_0p69 l=10
X235 dvdd.t199 a_35454_n291454.t41 por.t35 dvdd.t195 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X236 dvdd.t104 x2.Td_L.t8 x2.Td_Lb dvdd.t103 sky130_fd_pr__pfet_01v8 ad=0.217 pd=2.02 as=0.1155 ps=1.03 w=0.7 l=0.15
X237 a_28094_n290278.t5 x2.vbp1.t34 dvdd.t165 dvdd.t116 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X238 x1.VD.t2 x1.vo1.t2 x1.VY.t2 avss.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X239 a_28768_n287754# x2.Td_Sd.t12 dvdd.t76 dvdd.t75 sky130_fd_pr__pfet_01v8_hvt ad=0.196 pd=1.47 as=0.2352 ps=1.54 w=1.12 l=0.15
X240 a_18726_n286374# a_18492_n288774# dvss.t28 sky130_fd_pr__res_xhigh_po_0p69 l=10
X241 x2.x3.S1 x2.porbPre dvss.t389 dvss.t388 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
X242 a_29481_n287384# x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N dvdd.t161 dvdd.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.172775 ps=1.58 w=1 l=0.15
X243 a_35454_n291454.t5 a_35262_n291454.t13 dvss.t57 dvss.t56 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X244 a_28094_n290278.t4 x2.vbp1.t35 dvdd.t166 dvdd.t151 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X245 x2.Td_Sd.t3 a_25883_n288267.t7 dvss.t321 dvss.t320 sky130_fd_pr__nfet_01v8 ad=0.155 pd=1.62 as=0.0825 ps=0.83 w=0.5 l=0.15
X246 dvss.t421 a_30447_n287429# a_31115_n287366# dvss.t420 sky130_fd_pr__nfet_01v8 ad=0.126075 pd=1.1 as=0.15675 ps=1.67 w=0.55 l=0.15
X247 dvss.t11 x2.x3.S1B a_34073_n287091.t2 dvss.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=0.5
X248 x2.vbp1.t17 x2.vbp1.t16 dvdd.t272 dvdd.t33 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X249 dvdd.t133 a_28056_n288420# x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N dvdd.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X250 a_22237_n289908# a_22471_n292308# dvss.t140 sky130_fd_pr__res_xhigh_po_0p69 l=10
X251 a_30447_n287429# a_29688_n287709# a_30022_n287538# dvdd.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.22385 pd=1.7 as=0.39 ps=1.78 w=1 l=0.15
X252 dvdd.t80 a_35454_n291454.t42 por.t34 dvdd.t79 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X253 dvdd.t307 x2.porbPre a_35089_n289052# dvdd.t303 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.217 ps=2.02 w=0.7 l=0.15
X254 x2.VT3 dvss.t359 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X255 x2.Td_Lb x2.Td_L.t9 dvss.t110 dvss.t109 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.155 ps=1.62 w=0.5 l=0.15
X256 a_35454_n291454.t4 a_35262_n291454.t14 dvss.t59 dvss.t58 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X257 dvdd.t88 a_35469_n289052.t40 porb.t37 dvdd.t5 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X258 a_25216_n290828# a_24570_n290925.t4 x2.vbn1.t15 avdd.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
X259 dvss.t457 x2.VT2.t0 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X260 a_8822_n290308# avss.t14 avss.t13 sky130_fd_pr__res_xhigh_po_0p35 l=7
X261 dvss.t458 x2.VT3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X262 a_13030_n290763# x1.Vinp.t2 x1.VS avss.t65 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X263 porb_h[1].t26 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t25 avdd.t67 avdd.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X264 por.t10 a_35454_n291454.t43 dvss.t97 dvss.t96 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X265 a_20833_n289908# a_21067_n292308# dvss.t38 sky130_fd_pr__res_xhigh_po_0p69 l=10
X266 dvdd.t22 a_35277_n289052.t14 a_35469_n289052.t0 dvdd.t21 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X267 dvss.t1 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t26 porb_h[1].t11 dvss.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X268 x2.VT3 dvss.t358 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X269 dvss.t84 x2.Td_Sd.t13 a_29301_n287320# dvss.t83 sky130_fd_pr__nfet_01v8 ad=0.1212 pd=1.1 as=0.0504 ps=0.66 w=0.42 l=0.15
X270 a_30410_n291353# x2.VT2.t10 x2.VT3 dvss.t376 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.3
X271 a_28056_n288420# x2.delayPulse_digital_0/sky130_fd_sc_ls__xor2_1_0.X dvss.t289 dvss.t288 sky130_fd_pr__nfet_01v8 ad=0.1036 pd=1.02 as=0.12025 ps=1.065 w=0.74 l=0.15
X272 a_21534_n286374# a_21768_n288774# dvss.t29 sky130_fd_pr__res_xhigh_po_0p69 l=10
X273 dvss.t6 x2.Td_Sd.t14 a_28607_n287397# dvss.t5 sky130_fd_pr__nfet_01v8 ad=0.126075 pd=1.1 as=0.177375 ps=1.195 w=0.55 l=0.15
X274 dvss.t459 x2.VT3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X275 dvdd.t89 a_35469_n289052.t41 porb.t36 dvdd.t7 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X276 a_24270_n290121.t13 a_24270_n290121.t12 avdd.t98 avdd.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X277 dvss.t95 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t27 porb_h[0].t7 dvss.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X278 dvdd.t99 a_35469_n289052.t42 porb.t35 dvdd.t98 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X279 x2.Td_L.t4 a_32918_n290853.t5 dvdd.t18 dvdd.t17 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.217 ps=2.02 w=0.7 l=0.15
X280 a_9432_n286429# a_9598_n288829# avss.t34 sky130_fd_pr__res_xhigh_po_0p35 l=10
X281 por.t33 a_35454_n291454.t44 dvdd.t113 dvdd.t112 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X282 a_30728_n287754# a_29481_n287384# a_30447_n287429# dvdd.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.22385 ps=1.7 w=0.42 l=0.15
X283 dvss.t460 x2.VT3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X284 a_24270_n290121.t0 avdd.t25 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X285 avss.t50 x1.vo1.t3 a_9762_n292173# avss.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X286 avdd.t65 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t28 porb_h[1].t25 avdd.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X287 avdd.t3 a_34015_n286994.t5 a_34073_n287091.t1 avdd.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4205 pd=3.19 as=0.841 ps=6.38 w=2.9 l=0.5
X288 avdd.t63 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t29 porb_h[1].t24 avdd.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X289 avss.t8 x1.vbn.t1 x1.vbn.t2 avss.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X290 porb.t9 a_35469_n289052.t43 dvss.t105 dvss.t104 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X291 a_32918_n290853.t2 a_32248_n290278# dvdd.t178 dvdd.t176 sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.98 as=0.203 ps=1.98 w=0.7 l=0.15
X292 dvss.t461 x2.VT3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X293 a_19429_n289908# a_19195_n292308# dvss.t397 sky130_fd_pr__res_xhigh_po_0p69 l=10
X294 a_14804_n286429# a_14638_n288829# avss.t44 sky130_fd_pr__res_xhigh_po_0p35 l=10
X295 a_28868_n287397# x2.Td_L.t10 dvss.t281 dvss.t280 sky130_fd_pr__nfet_01v8 ad=0.0888 pd=0.98 as=0.126075 ps=1.1 w=0.74 l=0.15
X296 por.t9 a_35454_n291454.t45 dvss.t120 dvss.t119 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X297 a_21534_n286374# a_21300_n288774# dvss.t106 sky130_fd_pr__res_xhigh_po_0p69 l=10
X298 x2.VT2.t2 dvss.t332 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X299 a_5972_n290308.t4 a_5972_n290308.t3 avdd.t119 avdd.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X300 a_13808_n286429# a_13642_n288829# avss.t41 sky130_fd_pr__res_xhigh_po_0p35 l=10
X301 dvdd.t332 a_30447_n287429# a_31115_n287366# dvdd.t331 sky130_fd_pr__pfet_01v8_hvt ad=0.1862 pd=1.475 as=0.231 ps=2.23 w=0.84 l=0.15
X302 x2.VT3 dvss.t357 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X303 a_35469_n289052.t1 a_35277_n289052.t15 dvdd.t24 dvdd.t23 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X304 avdd.t85 a_24270_n290121.t10 a_24270_n290121.t11 avdd.t84 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X305 x1.vo1.t1 x1.vo.t3 w_15901_n291463# w_15901_n291463# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X306 a_36398_n287783.t2 x2.x3.aout.t4 avdd.t115 avdd.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3625 pd=2.79 as=0.725 ps=5.58 w=2.5 l=0.5
X307 porb.t34 a_35469_n289052.t44 dvdd.t291 dvdd.t96 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X308 a_25883_n288267.t0 dvss.t319 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X309 dvss.t462 x2.VT3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X310 x2.VT3 dvss.t356 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X311 dvdd.t202 x2.porPre a_35074_n291454# dvdd.t200 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.217 ps=2.02 w=0.7 l=0.15
X312 dvss.t425 x2.vbn1.t17 a_30410_n291353# dvss.t424 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.8
X313 avdd.t61 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t30 porb_h[0].t18 avdd.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X314 porb.t33 a_35469_n289052.t45 dvdd.t293 dvdd.t292 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X315 a_30031_n287373# a_29481_n287384# a_29895_n287373# dvss.t112 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1113 ps=0.95 w=0.42 l=0.15
X316 a_29671_n288104# a_29487_n288398# dvdd.t213 dvdd.t212 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.15 ps=1.3 w=1 l=0.15
X317 a_18961_n289908# a_18727_n292308# dvss.t316 sky130_fd_pr__res_xhigh_po_0p69 l=10
X318 a_21066_n286374# a_21300_n288774# dvss.t414 sky130_fd_pr__res_xhigh_po_0p69 l=10
X319 x2.VT2.t1 dvss.t417 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X320 dvss.t463 x2.VT3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X321 dvdd.t271 a_35454_n291454.t46 por.t32 dvdd.t270 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X322 x1.VS a_9762_n292173# x1.VY.t1 avss.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X323 dvss.t464 x2.VT2.t2 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X324 a_24253_n287224.t1 x2.din dvss.t429 dvss.t428 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.3
X325 a_30022_n287538# a_29895_n287373# dvdd.t286 dvdd.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=1.78 as=0.275 ps=2.55 w=1 l=0.15
X326 porb_h[0].t17 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t31 avdd.t60 avdd.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X327 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N a_28056_n288420# dvss.t150 dvss.t149 sky130_fd_pr__nfet_01v8 ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X328 a_25251_n288267.t0 dvss.t396 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X329 avdd.t122 a_24570_n290925.t0 sky130_fd_pr__cap_mim_m3_2 l=8 w=8
X330 x1.vo1.t0 x1.vo.t4 avss.t64 avss.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
X331 a_4566_n291516.t0 x1.vbn.t6 avss.t6 avss.t5 sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.3
X332 x1.VD.t8 x1.Vinn.t4 x1.VY.t6 avss.t69 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X333 dvdd.t249 x2.delayPulse_digital_0/sky130_fd_sc_ls__xor2_1_0.X a_28056_n288420# dvdd.t248 sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X334 a_13476_n286429# a_13642_n288829# avss.t28 sky130_fd_pr__res_xhigh_po_0p35 l=10
X335 x2.vbp1.t30 dvdd.t118 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X336 a_35454_n291454.t18 a_35262_n291454.t15 dvdd.t64 dvdd.t63 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X337 dvss.t8 x2.Td_Sd.t15 a_29487_n288398# dvss.t7 sky130_fd_pr__nfet_01v8 ad=0.162375 pd=1.255 as=0.2646 ps=2.4 w=0.74 l=0.15
X338 x1.Vinp.t0 a_12646_n288829# avss.t33 sky130_fd_pr__res_xhigh_po_0p35 l=10
X339 a_24570_n290925.t0 avdd.t99 sky130_fd_pr__cap_mim_m3_1 l=8 w=8
X340 a_35454_n291454.t17 a_35262_n291454.t16 dvdd.t236 dvdd.t90 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X341 dvss.t308 a_35454_n291454.t47 por.t8 dvss.t307 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X342 x1.VD.t0 a_9762_n292173# x1.VY.t0 avdd.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X343 dvdd.t16 a_30011_n288135# a_29966_n288037# dvdd.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.137125 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X344 avdd.t109 a_36398_n287783.t6 a_37002_n287783.t3 avdd.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.58 as=0.3625 ps=2.79 w=2.5 l=0.5
X345 a_22237_n289908# a_22003_n292308# dvss.t242 sky130_fd_pr__res_xhigh_po_0p69 l=10
X346 avdd.t59 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t32 porb_h[0].t21 avdd.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X347 a_35277_n289052.t0 a_35089_n289052# dvss.t213 dvss.t212 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X348 por.t31 a_35454_n291454.t48 dvdd.t69 dvdd.t53 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X349 dvss.t51 x2.x3.S1 a_34015_n286994.t0 dvss.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=0.5
X350 porb.t32 a_35469_n289052.t46 dvdd.t269 dvdd.t268 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X351 dvdd.t247 x2.delayPulse_digital_0/sky130_fd_sc_ls__xor2_1_0.X a_28056_n288420# dvdd.t246 sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X352 a_35454_n291454.t16 a_35262_n291454.t17 dvdd.t237 dvdd.t229 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X353 a_15914_n289870# x1.vo1.t4 avdd.t24 avdd.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X354 a_22938_n286374# a_22704_n288774# dvss.t157 sky130_fd_pr__res_xhigh_po_0p69 l=10
X355 x2.vbp1.t15 x2.vbp1.t14 dvdd.t267 dvdd.t144 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X356 avdd.t91 a_34073_n287091.t7 a_34015_n286994.t2 avdd.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4205 pd=3.19 as=0.841 ps=6.38 w=2.9 l=0.5
X357 porb.t8 a_35469_n289052.t47 dvss.t306 dvss.t305 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X358 por.t30 a_35454_n291454.t49 dvdd.t71 dvdd.t70 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X359 a_29895_n287373# a_29688_n287709# a_29214_n287320# dvss.t61 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=0.95 as=0.1113 ps=1.37 w=0.42 l=0.15
X360 dvdd.t218 x2.Td_Lb a_29211_n288416# dvdd.t217 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.05985 ps=0.705 w=0.42 l=0.15
X361 dvdd.t288 x2.VT2.t11 x2.VT3 dvdd.t287 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X362 a_25883_n288267.t2 a_25567_n288267.t5 dvss.t3 dvss.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
X363 a_30814_n289746# a_24253_n287224.t7 x2.VT2.t5 dvdd.t317 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X364 a_21769_n289908# a_22003_n292308# dvss.t179 sky130_fd_pr__res_xhigh_po_0p69 l=10
X365 a_9100_n286429# a_8934_n288829# avss.t21 sky130_fd_pr__res_xhigh_po_0p35 l=10
X366 a_35469_n289052.t12 a_35277_n289052.t16 dvdd.t206 dvdd.t205 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X367 porb_h[0].t20 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t33 avdd.t58 avdd.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X368 dvss.t373 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t34 porb_h[1].t10 dvss.t372 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X369 a_8104_n286429# a_7938_n288829# avss.t70 sky130_fd_pr__res_xhigh_po_0p35 l=10
X370 por.t29 a_35454_n291454.t50 dvdd.t333 dvdd.t295 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X371 a_20365_n289908# a_20599_n292308# dvss.t118 sky130_fd_pr__res_xhigh_po_0p69 l=10
X372 a_22470_n286374# a_22704_n288774# dvss.t124 sky130_fd_pr__res_xhigh_po_0p69 l=10
X373 dvdd.t241 x2.Td_L.t11 a_28768_n287754# dvdd.t240 sky130_fd_pr__pfet_01v8_hvt ad=0.2352 pd=1.54 as=0.3752 ps=2.91 w=1.12 l=0.15
X374 a_13030_n290763# x1.Vinp.t3 x1.VS avss.t65 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X375 a_29298_n288416# x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtp_1_0.D a_29211_n288416# dvss.t413 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X376 dvss.t209 x2.vbn1.t7 x2.vbn1.t8 dvss.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.8
X377 dvdd.t74 a_35469_n289052.t48 porb.t31 dvdd.t73 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X378 dvss.t241 a_35277_n289052.t17 a_35469_n289052.t13 dvss.t240 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X379 a_30779_n287655# x2.Td_Sd.t16 dvdd.t10 dvdd.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0819 ps=0.81 w=0.42 l=0.15
X380 x2.porbPre a_31115_n287366# dvdd.t142 dvdd.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.3192 pd=2.81 as=0.1862 ps=1.475 w=1.12 l=0.15
X381 a_30022_n287538# a_29895_n287373# dvss.t341 dvss.t340 sky130_fd_pr__nfet_01v8 ad=0.1073 pd=1.03 as=0.240325 ps=1.715 w=0.74 l=0.15
X382 por.t28 a_35454_n291454.t51 dvdd.t334 dvdd.t148 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X383 dvdd.t238 a_35262_n291454.t18 a_35454_n291454.t15 dvdd.t94 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X384 x2.vbp1.t13 x2.vbp1.t12 dvdd.t117 dvdd.t116 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X385 a_7996_n292010# x1.vbn.t7 a_5972_n290308.t1 avss.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X386 x2.VT2.t2 dvss.t331 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X387 a_20365_n289908# a_20131_n292308# dvss.t39 sky130_fd_pr__res_xhigh_po_0p69 l=10
X388 x2.vbp1.t11 x2.vbp1.t10 dvdd.t152 dvdd.t151 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X389 a_36398_n287783.t3 x2.x3.aout.t5 dvss.t411 dvss.t410 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X390 dvdd.t298 x2.vbp1.t36 a_28094_n290278.t3 dvdd.t55 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X391 dvss.t287 x2.delayPulse_digital_0/sky130_fd_sc_ls__xor2_1_0.X a_28056_n288420# dvss.t286 sky130_fd_pr__nfet_01v8 ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X392 dvss.t393 a_35277_n289052.t18 a_35469_n289052.t16 dvss.t392 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X393 porb_h[0].t6 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t35 dvss.t375 dvss.t374 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X394 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N a_28056_n288420# dvdd.t131 dvdd.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X395 a_30447_n288420# a_29671_n288104# a_30011_n288135# dvss.t263 sky130_fd_pr__nfet_01v8 ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X396 dvss.t337 a_35074_n291454# a_35262_n291454.t1 dvss.t336 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X397 a_15914_n289870# x1.vo1.t5 avss.t37 avss.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X398 dvss.t251 a_27214_n288191# a_27214_n288191# dvss.t250 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
X399 a_30657_n288413# a_29487_n288398# a_30447_n288420# dvss.t255 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X400 x2.VT2.t1 dvss.t416 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X401 dvdd.t282 a_35074_n291454# a_35262_n291454.t3 dvdd.t280 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X402 dvss.t80 a_35469_n289052.t49 porb.t7 dvss.t79 sky130_fd_pr__nfet_01v8 ad=0.155 pd=1.62 as=0.0825 ps=0.83 w=0.5 l=0.15
X403 dvss.t406 a_35454_n291454.t52 por.t7 dvss.t405 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X404 dvdd.t20 a_32918_n290853.t6 x2.Td_L.t3 dvdd.t19 sky130_fd_pr__pfet_01v8 ad=0.217 pd=2.02 as=0.1155 ps=1.03 w=0.7 l=0.15
X405 a_19897_n289908# a_20131_n292308# dvss.t174 sky130_fd_pr__res_xhigh_po_0p69 l=10
X406 a_35277_n289052.t3 a_35089_n289052# dvdd.t189 dvdd.t188 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X407 dvss.t129 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t36 porb_h[1].t9 dvss.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X408 a_18493_n289908# a_18727_n292308# dvss.t123 sky130_fd_pr__res_xhigh_po_0p69 l=10
X409 a_14472_n286429# a_14638_n288829# avss.t47 sky130_fd_pr__res_xhigh_po_0p35 l=10
X410 dvdd.t319 a_35454_n291454.t53 por.t27 dvdd.t259 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X411 a_20598_n286374# a_20832_n288774# dvss.t400 sky130_fd_pr__res_xhigh_po_0p69 l=10
X412 a_25567_n288267.t1 a_25251_n288267.t6 dvss.t395 dvss.t394 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
X413 x1.vbn.t0 a_5972_n290308.t5 avdd.t117 avdd.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X414 a_30075_n288356# a_30011_n288135# a_29997_n288356# dvss.t18 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X415 porb.t30 a_35469_n289052.t50 dvdd.t183 dvdd.t162 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X416 dvss.t137 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t37 porb_h[0].t5 dvss.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X417 dvdd.t197 a_35454_n291454.t54 por.t26 dvdd.t79 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X418 x2.VT3 dvss.t355 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X419 a_30011_n288135# a_29876_n288037# dvdd.t339 dvdd.t338 sky130_fd_pr__pfet_01v8_hvt ad=0.190625 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X420 dvdd.t300 x2.vbp1.t37 a_28094_n290278.t2 dvdd.t299 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X421 avdd.t57 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t38 porb_h[0].t19 avdd.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X422 dvss.t211 a_35469_n289052.t51 porb.t6 dvss.t210 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X423 x2.Td_L.t0 a_32918_n290853.t7 dvss.t206 dvss.t205 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.155 ps=1.62 w=0.5 l=0.15
X424 dvss.t465 x2.VT3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X425 dvss.t268 a_35262_n291454.t19 a_35454_n291454.t3 dvss.t267 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X426 dvdd.t198 a_35454_n291454.t55 por.t25 dvdd.t146 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X427 x1.VD.t7 x1.Vinn.t5 x1.VY.t5 avss.t69 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X428 dvdd.t187 a_35089_n289052# a_35277_n289052.t2 dvdd.t186 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X429 x2.vbp1.t29 x2.vbp2 x2.vbp2 dvdd.t13 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X430 x2.Td_S.t3 a_24253_n287224.t8 dvdd.t316 dvdd.t174 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X431 x2.VT3 dvss.t354 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X432 dvdd.t312 a_35277_n289052.t19 a_35469_n289052.t17 dvdd.t311 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X433 dvss.t466 x2.VT3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X434 w_15901_n291463# w_15901_n291463# avdd.t27 avdd.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X435 dvss.t285 x2.delayPulse_digital_0/sky130_fd_sc_ls__xor2_1_0.X a_28056_n288420# dvss.t284 sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.065 as=0.2109 ps=2.05 w=0.74 l=0.15
X436 a_35454_n291454.t2 a_35262_n291454.t20 dvss.t270 dvss.t269 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X437 dvss.t467 a_25883_n288267.t0 sky130_fd_pr__cap_mim_m3_2 l=10 w=10
X438 dvdd.t264 a_35469_n289052.t52 porb.t29 dvdd.t31 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X439 avdd.t87 a_24270_n290121.t8 a_24270_n290121.t9 avdd.t86 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X440 a_30447_n288420# a_29487_n288398# a_30011_n288135# dvdd.t211 sky130_fd_pr__pfet_01v8_hvt ad=0.23015 pd=1.73 as=0.190625 ps=1.505 w=1 l=0.15
X441 dvss.t468 x2.VT2.t3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X442 a_21769_n289908# a_21535_n292308# dvss.t72 sky130_fd_pr__res_xhigh_po_0p69 l=10
X443 a_14472_n286429# a_14306_n288829# avss.t12 sky130_fd_pr__res_xhigh_po_0p35 l=10
X444 a_30699_n288291# x2.Td_Lb dvdd.t216 dvdd.t215 sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X445 a_35454_n291454.t14 a_35262_n291454.t21 dvdd.t225 dvdd.t224 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X446 a_13476_n286429# a_13310_n288829# avss.t71 sky130_fd_pr__res_xhigh_po_0p35 l=10
X447 dvdd.t314 a_35277_n289052.t20 a_35469_n289052.t18 dvdd.t192 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X448 a_24253_n287224.t3 x2.din dvdd.t337 dvdd.t335 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X449 dvss.t148 a_28056_n288420# x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N dvss.t147 sky130_fd_pr__nfet_01v8 ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X450 dvdd.t266 a_35469_n289052.t53 porb.t28 dvdd.t265 sky130_fd_pr__pfet_01v8 ad=0.217 pd=2.02 as=0.1155 ps=1.03 w=0.7 l=0.15
X451 dvss.t116 x2.vbn1.t5 x2.vbn1.t6 dvss.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X452 dvss.t469 x2.VT3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X453 avdd.t56 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t39 porb_h[1].t23 avdd.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X454 a_25251_n288267.t2 x2.Td_S.t5 dvss.t45 dvss.t44 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
X455 a_21301_n289908# a_21535_n292308# dvss.t34 sky130_fd_pr__res_xhigh_po_0p69 l=10
X456 x2.din a_15914_n289870# avss.t67 avss.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X457 x2.Td_S.t0 a_24253_n287224.t9 dvss.t399 dvss.t398 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.3
X458 a_29671_n288104# a_29487_n288398# dvss.t254 dvss.t253 sky130_fd_pr__nfet_01v8 ad=0.2183 pd=2.07 as=0.162375 ps=1.255 w=0.74 l=0.15
X459 porb_h[1].t8 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t40 dvss.t93 dvss.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X460 x1.VS x1.vo1.t6 x1.VY.t3 avdd.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X461 porb.t5 a_35469_n289052.t54 dvss.t192 dvss.t191 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X462 a_29688_n287709# a_29481_n287384# dvdd.t109 dvdd.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.40345 pd=2.86 as=0.295 ps=2.59 w=1 l=0.15
X463 dvss.t470 x2.VT3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X464 dvdd.t201 x2.porPre a_35074_n291454# dvdd.t200 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.217 ps=2.02 w=0.7 l=0.15
X465 por.t6 a_35454_n291454.t56 dvss.t404 dvss.t403 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X466 a_11424_n286429# a_11258_n288829# avss.t16 sky130_fd_pr__res_xhigh_po_0p35 l=10
X467 x2.x3.S1B x2.x3.S1 dvdd.t60 dvdd.t59 sky130_fd_pr__pfet_01v8 ad=0.217 pd=2.02 as=0.1155 ps=1.03 w=0.7 l=0.15
X468 dvss.t323 a_25883_n288267.t8 x2.Td_Sd.t4 dvss.t322 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.155 ps=1.62 w=0.5 l=0.15
X469 x2.VT3 dvss.t353 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X470 a_35469_n289052.t19 a_35277_n289052.t21 dvdd.t315 dvdd.t27 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X471 a_10428_n286429# a_10262_n288829# avss.t40 sky130_fd_pr__res_xhigh_po_0p35 l=10
X472 x2.vbn1.t4 x2.vbn1.t3 dvss.t20 dvss.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X473 a_21301_n289908# a_21067_n292308# dvss.t27 sky130_fd_pr__res_xhigh_po_0p69 l=10
X474 porb_h[1].t22 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t41 avdd.t54 avdd.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X475 dvdd.t318 a_35454_n291454.t57 por.t24 dvdd.t270 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X476 x2.Td_S.t2 a_24253_n287224.t10 dvdd.t175 dvdd.t174 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X477 a_30699_n288291# a_30447_n288420# a_30837_n288413# dvss.t290 sky130_fd_pr__nfet_01v8 ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X478 dvdd.t168 a_35469_n289052.t55 porb.t27 dvdd.t29 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X479 x2.VT3 dvss.t352 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X480 dvss.t312 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t42 porb_h[1].t7 dvss.t311 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X481 dvss.t471 x2.VT2.t1 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X482 dvss.t272 a_35262_n291454.t22 a_35454_n291454.t1 dvss.t271 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X483 dvss.t472 x2.VT2.t2 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X484 a_32248_n290278# x2.VT3 dvss.t351 dvss.t350 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.3
X485 dvss.t314 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t43 porb_h[0].t4 dvss.t313 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X486 a_28056_n288420# x2.delayPulse_digital_0/sky130_fd_sc_ls__xor2_1_0.X dvdd.t245 dvdd.t244 sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X487 a_24253_n287224.t2 x2.din dvdd.t336 dvdd.t335 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X488 dvss.t165 a_35454_n291454.t58 por.t5 dvss.t164 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X489 a_35454_n291454.t13 a_35262_n291454.t23 dvdd.t226 dvdd.t63 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X490 avdd.t15 x1.vo1.t7 a_9762_n292173# avdd.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X491 dvdd.t204 a_30022_n287538# a_29998_n287709# dvdd.t203 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0504 ps=0.66 w=0.42 l=0.15
X492 a_35469_n289052.t14 a_35277_n289052.t22 dvdd.t310 dvdd.t25 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X493 avdd.t52 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t44 porb_h[1].t21 avdd.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X494 dvss.t473 x2.VT2.t2 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X495 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t2 a_37002_n287783.t5 avdd.t105 avdd.t104 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3625 pd=2.79 as=0.725 ps=5.58 w=2.5 l=0.5
X496 dvss.t159 a_34073_n287091.t8 x2.x3.aout.t0 dvss.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=0.5
X497 porb_h[1].t6 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t45 dvss.t55 dvss.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X498 a_28094_n290278.t1 x2.vbp1.t38 dvdd.t41 dvdd.t40 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X499 porb.t26 a_35469_n289052.t56 dvdd.t101 dvdd.t100 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X500 porb.t25 a_35469_n289052.t57 dvdd.t102 dvdd.t38 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X501 a_8436_n286429# a_8602_n288829# avss.t17 sky130_fd_pr__res_xhigh_po_0p35 l=10
X502 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N a_28056_n288420# dvdd.t129 dvdd.t128 sky130_fd_pr__pfet_01v8_hvt ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X503 a_10096_n286429# a_10262_n288829# avss.t26 sky130_fd_pr__res_xhigh_po_0p35 l=10
X504 avss.t73 a_7606_n288829# avss.t72 sky130_fd_pr__res_xhigh_po_0p35 l=10
X505 dvdd.t208 a_27214_n288191# x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtp_1_0.D dvdd.t207 sky130_fd_pr__pfet_01v8 ad=0.155 pd=1.62 as=0.0825 ps=0.83 w=0.5 l=0.15
X506 dvdd.t228 a_35262_n291454.t24 a_35454_n291454.t12 dvdd.t227 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X507 a_35454_n291454.t11 a_35262_n291454.t25 dvdd.t230 dvdd.t229 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X508 avdd.t50 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t46 porb_h[0].t16 avdd.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X509 a_22705_n289908# a_22939_n292308# dvss.t239 sky130_fd_pr__res_xhigh_po_0p69 l=10
X510 dvdd.t105 x2.Td_L.t12 x2.Td_Lb dvdd.t103 sky130_fd_pr__pfet_01v8 ad=0.217 pd=2.02 as=0.1155 ps=1.03 w=0.7 l=0.15
X511 porb_h[1].t20 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t47 avdd.t49 avdd.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X512 dvdd.t306 x2.porbPre x2.x3.S1 dvdd.t305 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.217 ps=2.02 w=0.7 l=0.15
X513 x2.VT3 dvss.t349 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X514 x2.VT2.t0 dvss.t196 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X515 x2.VT3 dvss.t348 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X516 por.t23 a_35454_n291454.t59 dvdd.t153 dvdd.t70 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X517 a_35469_n289052.t15 a_35277_n289052.t23 dvss.t391 dvss.t390 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X518 porb.t24 a_35469_n289052.t58 dvdd.t87 dvdd.t45 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X519 a_13449_n292106.t0 avdd.t123 a_13030_n290763# avss.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
X520 x2.VT3 dvss.t347 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X521 avdd.t12 x1.vo1.t8 a_15914_n289870# avdd.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X522 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t0 a_37002_n287783.t6 dvss.t31 dvss.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X523 porb.t4 a_35469_n289052.t59 dvss.t101 dvss.t100 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X524 dvdd.t56 x2.vbp1.t8 x2.vbp1.t9 dvdd.t55 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X525 a_22705_n289908# a_22471_n292308# dvss.t238 sky130_fd_pr__res_xhigh_po_0p69 l=10
X526 porb_h[0].t25 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t48 avdd.t47 avdd.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X527 porb_h[0].t24 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t49 avdd.t46 avdd.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X528 a_30779_n287655# a_30447_n287429# a_30917_n287365# dvss.t419 sky130_fd_pr__nfet_01v8 ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X529 x2.VT2.t3 dvss.t327 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X530 porb.t23 a_35469_n289052.t60 dvdd.t58 dvdd.t57 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X531 dvdd.t330 a_30447_n287429# a_30779_n287655# dvdd.t329 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0.063 ps=0.72 w=0.42 l=0.15
X532 dvss.t474 a_25251_n288267.t0 sky130_fd_pr__cap_mim_m3_2 l=10 w=10
X533 dvdd.t78 a_35277_n289052.t24 a_35469_n289052.t4 dvdd.t77 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X534 a_24270_n290121.t7 a_24270_n290121.t6 avdd.t29 avdd.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.8
X535 x2.VT2.t0 dvss.t195 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X536 por.t22 a_35454_n291454.t60 dvdd.t149 dvdd.t148 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X537 x2.Td_Lb x2.Td_L.t13 dvdd.t107 dvdd.t106 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.217 ps=2.02 w=0.7 l=0.15
X538 x2.Td_Sd.t5 a_25883_n288267.t9 dvdd.t278 dvdd.t273 sky130_fd_pr__pfet_01v8 ad=0.217 pd=2.02 as=0.1155 ps=1.03 w=0.7 l=0.15
X539 a_29214_n287320# x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtp_1_0.D dvdd.t326 dvdd.t325 sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.1218 ps=1.42 w=0.42 l=0.15
X540 dvss.t47 a_35469_n289052.t61 porb.t3 dvss.t46 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X541 dvss.t475 x2.VT3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X542 a_19194_n286374# a_18960_n288774# dvss.t262 sky130_fd_pr__res_xhigh_po_0p69 l=10
X543 dvdd.t127 a_28056_n288420# x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N dvdd.t126 sky130_fd_pr__pfet_01v8_hvt ad=0.1876 pd=1.455 as=0.168 ps=1.42 w=1.12 l=0.15
X544 avdd.t93 a_24270_n290121.t18 a_25216_n290828# avdd.t92 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
X545 dvss.t476 x2.VT2.t0 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X546 por.t21 a_35454_n291454.t61 dvdd.t150 dvdd.t82 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X547 x2.VT2.t3 dvss.t326 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X548 dvdd.t302 x2.vbp1.t6 x2.vbp1.t7 dvdd.t299 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X549 avdd.t22 a_34073_n287091.t9 x2.x3.aout.t1 avdd.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4205 pd=3.19 as=0.841 ps=6.38 w=2.9 l=0.5
X550 a_4566_n290308.t2 a_4566_n290308.t1 avdd.t110 avdd.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X551 dvss.t477 x2.VT2.t0 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X552 dvdd.t281 a_35074_n291454# a_35262_n291454.t2 dvdd.t280 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X553 a_29876_n288037# a_29671_n288104# a_29211_n288416# dvdd.t222 sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.1218 ps=1.42 w=0.42 l=0.15
X554 dvss.t91 a_35277_n289052.t25 a_35469_n289052.t5 dvss.t90 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X555 x2.VT2.t0 dvss.t194 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X556 a_28607_n287397# x2.Td_L.t14 dvss.t369 dvss.t368 sky130_fd_pr__nfet_01v8 ad=0.177375 pd=1.195 as=0.33275 ps=2.31 w=0.55 l=0.15
X557 dvdd.t125 a_28056_n288420# x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N dvdd.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.3304 pd=2.83 as=0.1764 ps=1.435 w=1.12 l=0.15
X558 a_31045_n288085# a_30447_n288420# dvdd.t253 dvdd.t252 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X559 a_32918_n290853.t1 a_32248_n290278# dvdd.t177 dvdd.t176 sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.98 as=0.203 ps=1.98 w=0.7 l=0.15
X560 w_31992_n290497# x2.vbp2 a_28094_n290278.t8 dvdd.t12 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X561 a_30112_n289746# x2.vbp1.t39 dvdd.t42 dvdd.t13 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X562 a_37002_n287783.t2 a_36398_n287783.t7 avdd.t107 avdd.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3625 pd=2.79 as=0.725 ps=5.58 w=2.5 l=0.5
X563 x2.din a_15914_n289870# dvdd.t322 dvdd.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X564 dvss.t387 x2.porbPre a_35089_n289052# dvss.t386 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.155 ps=1.62 w=0.5 l=0.15
X565 dvdd.t260 a_35454_n291454.t62 por.t20 dvdd.t259 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X566 a_20833_n289908# a_20599_n292308# dvss.t432 sky130_fd_pr__res_xhigh_po_0p69 l=10
X567 avdd.t45 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t50 porb_h[1].t19 avdd.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X568 dvdd.t232 a_35262_n291454.t26 a_35454_n291454.t10 dvdd.t231 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X569 x2.vbp2 x2.vbp2 x2.vbp1.t28 dvdd.t11 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X570 avdd.t17 avdd.t16 a_14970_n288829# avss.t15 sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.9
X571 x2.VT2.t4 a_24253_n287224.t11 dvss.t202 dvss.t201 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.3
X572 dvss.t186 a_35469_n289052.t62 porb.t2 dvss.t185 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X573 avdd.t7 a_24270_n290121.t4 a_24270_n290121.t5 avdd.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.8
X574 x2.VT2.t3 dvss.t325 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X575 dvss.t310 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t51 porb_h[0].t3 dvss.t309 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X576 a_14804_n286429# a_14970_n288829# avss.t46 sky130_fd_pr__res_xhigh_po_0p35 l=10
X577 dvdd.t261 a_35454_n291454.t63 por.t19 dvdd.t255 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X578 a_11092_n286429# a_11258_n288829# avss.t29 sky130_fd_pr__res_xhigh_po_0p35 l=10
X579 dvss.t283 a_31045_n288085# x2.porPre dvss.t282 sky130_fd_pr__nfet_01v8 ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X580 avss.t4 x1.vbn.t8 x1.VS avss.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X581 a_13808_n286429# a_13974_n288829# avss.t74 sky130_fd_pr__res_xhigh_po_0p35 l=10
X582 dvdd.t147 a_35454_n291454.t64 por.t18 dvdd.t146 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X583 x2.VT2.t0 dvss.t193 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X584 a_12812_n286429# a_12978_n288829# avss.t45 sky130_fd_pr__res_xhigh_po_0p35 l=10
X585 porb_h[1].t5 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t52 dvss.t217 dvss.t216 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X586 porb_h[1].t4 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t53 dvss.t219 dvss.t218 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X587 dvss.t478 x2.VT3 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X588 x2.delayPulse_digital_0/sky130_fd_sc_ls__xor2_1_0.X x2.Td_Sd.t17 a_28868_n287397# dvss.t37 sky130_fd_pr__nfet_01v8 ad=0.1554 pd=1.16 as=0.0888 ps=0.98 w=0.74 l=0.15
X589 a_29301_n287320# x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtp_1_0.D a_29214_n287320# dvss.t412 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X590 dvss.t146 a_28056_n288420# x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N dvss.t145 sky130_fd_pr__nfet_01v8 ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X591 dvss.t188 a_35469_n289052.t63 porb.t1 dvss.t187 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X592 a_30731_n287365# a_29688_n287709# a_30447_n287429# dvss.t60 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.3067 ps=2.01 w=0.42 l=0.15
X593 dvss.t163 a_35454_n291454.t65 por.t4 dvss.t162 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X594 dvdd.t251 a_30447_n288420# a_30699_n288291# dvdd.t250 sky130_fd_pr__pfet_01v8_hvt ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X595 x2.VT2.t3 dvss.t324 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X596 x1.vo.t5 x1.vt.t1 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X597 dvdd.t173 a_35277_n289052.t26 a_35469_n289052.t6 dvdd.t21 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X598 dvdd.t158 a_35469_n289052.t64 porb.t22 dvdd.t47 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X599 a_8822_n290308# a_8656_n292108# avss.t35 sky130_fd_pr__res_xhigh_po_0p35 l=7
X600 a_4566_n291516.t2 a_4566_n291516.t1 a_4508_n291419.t2 avdd.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X601 dvdd.t85 a_35454_n291454.t66 por.t17 dvdd.t84 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X602 a_35454_n291454.t9 a_35262_n291454.t27 dvdd.t233 dvdd.t224 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X603 a_32248_n290278# x2.VT3 w_31992_n290497# w_31992_n290497# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X604 porb_h[0].t23 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t54 avdd.t43 avdd.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X605 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N a_28056_n288420# dvss.t144 dvss.t143 sky130_fd_pr__nfet_01v8 ad=0.10545 pd=1.025 as=0.1554 ps=1.16 w=0.74 l=0.15
X606 porb_h[0].t31 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t55 avdd.t41 avdd.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X607 dvdd.t159 a_35469_n289052.t65 porb.t21 dvdd.t98 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X608 x2.x3.S1B x2.x3.S1 dvss.t49 dvss.t48 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
X609 a_10760_n286429# a_10926_n288829# avss.t38 sky130_fd_pr__res_xhigh_po_0p35 l=10
X610 dvss.t244 x2.x3.aout.t6 a_36398_n287783.t1 dvss.t243 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X611 x2.VT3 dvss.t346 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X612 a_35469_n289052.t7 a_35277_n289052.t27 dvss.t200 dvss.t199 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X613 a_9432_n286429# a_9266_n288829# avss.t51 sky130_fd_pr__res_xhigh_po_0p35 l=10
X614 a_35262_n291454.t0 a_35074_n291454# dvss.t335 dvss.t334 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X615 a_11092_n286429# a_10926_n288829# avss.t75 sky130_fd_pr__res_xhigh_po_0p35 l=10
X616 dvdd.t349 x2.vbp1.t30 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X617 a_8436_n286429# a_8270_n288829# avss.t23 sky130_fd_pr__res_xhigh_po_0p35 l=10
X618 x2.VT2.t2 dvss.t330 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X619 dvss.t24 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t56 porb_h[0].t2 dvss.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X620 a_10096_n286429# a_9930_n288829# avss.t42 sky130_fd_pr__res_xhigh_po_0p35 l=10
X621 porb.t0 a_35469_n289052.t66 dvss.t103 dvss.t102 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X622 dvss.t182 dvdd.t350 dvss.t181 dvss.t180 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0 ps=0 w=0.42 l=1
X623 por.t3 a_35454_n291454.t67 dvss.t99 dvss.t98 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X624 dvdd.t304 x2.porbPre a_35089_n289052# dvdd.t303 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.217 ps=2.02 w=0.7 l=0.15
X625 dvss.t479 x2.vbn1.t0 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X626 porb.t20 a_35469_n289052.t67 dvdd.t97 dvdd.t96 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X627 avdd.t39 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t57 porb_h[0].t30 avdd.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X628 dvss.t480 a_25567_n288267.t0 sky130_fd_pr__cap_mim_m3_2 l=10 w=10
X629 dvdd.t68 a_30699_n288291# a_30649_n288001# dvdd.t67 sky130_fd_pr__pfet_01v8_hvt ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X630 x2.VT2.t1 dvss.t415 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X631 x2.VT3 dvss.t345 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X632 dvdd.t6 a_35469_n289052.t68 porb.t19 dvdd.t5 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X633 a_7996_n292010# x1.vbn.t9 a_5972_n290308.t0 avss.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X634 por.t2 a_35454_n291454.t68 dvss.t385 dvss.t384 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X635 x2.vbp2 x2.vbn1.t18 dvss.t378 dvss.t377 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
X636 x2.vbp1.t5 x2.vbp1.t4 dvdd.t86 dvdd.t40 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X637 dvdd.t2 dvss.t481 dvdd.t1 dvdd.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=1
X638 avdd.t10 a_13449_n292106.t1 a_13449_n292106.t2 avdd.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
X639 a_10760_n286429# a_10594_n288829# avss.t43 sky130_fd_pr__res_xhigh_po_0p35 l=10
X640 dvdd.t123 a_28056_n288420# x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N dvdd.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X641 a_29876_n288037# a_29487_n288398# a_29211_n288416# dvss.t252 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X642 por.t16 a_35454_n291454.t69 dvdd.t301 dvdd.t257 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X643 porb_h[0].t29 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t58 avdd.t37 avdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X644 dvss.t22 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t59 porb_h[1].t3 dvss.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.2025 pd=2.04 as=0.105 ps=1.03 w=0.75 l=0.5
X645 dvdd.t8 a_35469_n289052.t69 porb.t18 dvdd.t7 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X646 avss.t2 x1.vbn.t10 x1.VS avss.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X647 x2.VT3 dvss.t344 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X648 a_8104_n286429# a_8270_n288829# avss.t56 sky130_fd_pr__res_xhigh_po_0p35 l=10
X649 a_23173_n289908# vbg.t0 a_24570_n290925.t1 dvss.t237 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X650 a_25883_n288267.t3 a_25567_n288267.t6 dvdd.t221 dvdd.t3 sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.98 as=0.203 ps=1.98 w=0.7 l=0.15
X651 dvss.t371 x2.Td_L.t15 x2.Td_Lb dvss.t370 sky130_fd_pr__nfet_01v8 ad=0.155 pd=1.62 as=0.0825 ps=0.83 w=0.5 l=0.15
X652 dvss.t274 a_35262_n291454.t28 a_35454_n291454.t0 dvss.t273 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X653 avdd.t101 a_24270_n290121.t2 a_24270_n290121.t3 avdd.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X654 dvss.t482 x2.VT2.t1 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X655 a_18258_n286374# a_18492_n288774# dvss.t383 sky130_fd_pr__res_xhigh_po_0p69 l=10
X656 dvdd.t254 x2.vbp1.t2 x2.vbp1.t3 dvdd.t156 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X657 x1.vt.t0 avdd.t124 x1.VD.t1 avss.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
X658 avdd.t35 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t60 porb_h[1].t18 avdd.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X659 a_30447_n287429# a_29481_n287384# a_30022_n287538# dvss.t111 sky130_fd_pr__nfet_01v8 ad=0.3067 pd=2.01 as=0.1073 ps=1.03 w=0.74 l=0.15
X660 dvss.t380 x2.vbn1.t19 a_30410_n291353# dvss.t379 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X661 porb_h[1].t2 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t61 dvss.t266 dvss.t265 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X662 porb_h[1].t1 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t62 dvss.t133 dvss.t132 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X663 dvdd.t263 x2.vbp1.t0 x2.vbp1.t1 dvdd.t262 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X664 dvss.t298 a_35454_n291454.t70 por.t1 dvss.t297 sky130_fd_pr__nfet_01v8 ad=0.155 pd=1.62 as=0.0825 ps=0.83 w=0.5 l=0.15
X665 a_35469_n289052.t10 a_35277_n289052.t28 dvdd.t194 dvdd.t23 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X666 dvss.t483 x2.VT2.t1 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X667 dvdd.t234 a_35262_n291454.t29 a_35454_n291454.t8 dvdd.t227 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X668 a_22938_n286374# dvss.t246 dvss.t245 sky130_fd_pr__res_xhigh_po_0p69 l=10
X669 dvss.t142 a_28056_n288420# x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N dvss.t141 sky130_fd_pr__nfet_01v8 ad=0.2627 pd=2.19 as=0.10545 ps=1.025 w=0.74 l=0.15
X670 dvss.t257 x2.Td_Lb a_29298_n288416# dvss.t256 sky130_fd_pr__nfet_01v8 ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X671 a_25251_n288267.t3 x2.Td_S.t6 dvdd.t313 dvdd.t49 sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.98 as=0.203 ps=1.98 w=0.7 l=0.15
X672 porb_h[0].t1 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t63 dvss.t135 dvss.t134 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X673 avdd.t103 a_37002_n287783.t7 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t3 avdd.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.58 as=0.3625 ps=2.79 w=2.5 l=0.5
X674 dvss.t127 a_30779_n287655# a_30731_n287365# dvss.t126 sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.0504 ps=0.66 w=0.42 l=0.15
X675 a_35469_n289052.t11 a_35277_n289052.t29 dvss.t227 dvss.t226 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X676 porb.t17 a_35469_n289052.t70 dvdd.t343 dvdd.t268 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X677 dvdd.t179 a_32918_n290853.t8 x2.Td_L.t2 dvdd.t19 sky130_fd_pr__pfet_01v8 ad=0.217 pd=2.02 as=0.1155 ps=1.03 w=0.7 l=0.15
X678 porb.t16 a_35469_n289052.t71 dvdd.t344 dvdd.t292 sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X679 porb_h[1].t17 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t64 avdd.t33 avdd.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X680 a_30410_n291353# x2.vbn1.t20 dvss.t89 dvss.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X681 porb_h[1].t16 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t65 avdd.t31 avdd.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X682 x1.VD.t3 x1.Vinn.t6 x1.VS avss.t19 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X683 x1.VD.t6 x1.Vinn.t7 x1.VY.t4 avss.t20 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X684 dvss.t131 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t66 porb_h[1].t0 dvss.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X685 dvss.t300 a_35454_n291454.t71 por.t0 dvss.t299 sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X686 x2.VT3 dvss.t343 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X687 dvss.t484 x2.VT2.t0 sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X688 x2.vbn1.t2 x2.vbn1.t1 dvss.t172 dvss.t171 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X689 dvdd.t185 x2.vbp1.t40 a_28094_n290278.t0 dvdd.t184 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X690 dvss.t87 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t67 porb_h[0].t0 dvss.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X691 dvss.t427 x2.din a_24253_n287224.t0 dvss.t426 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.3
X692 dvss.t74 a_30699_n288291# a_30657_n288413# dvss.t73 sky130_fd_pr__nfet_01v8 ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
R0 dvss.n1038 dvss.n1037 205907
R1 dvss.t350 dvss.n754 164476
R2 dvss.n1278 dvss.n1257 126229
R3 dvss.n1278 dvss.n1258 120611
R4 dvss.n1311 dvss.n47 93411
R5 dvss.n1274 dvss.n1258 93404.6
R6 dvss.n1038 dvss.n1035 90168.1
R7 dvss.n1274 dvss.n1261 77113.4
R8 dvss.n1265 dvss.n1257 54654.1
R9 dvss.n1414 dvss.n25 42361.3
R10 dvss.n507 dvss.n458 40791.1
R11 dvss.n1314 dvss.n1311 37112.5
R12 dvss.n1062 dvss.n1061 33058.4
R13 dvss.n1265 dvss.n1261 32711.6
R14 dvss.n1277 dvss.n1259 29011.1
R15 dvss.n1161 dvss.n786 25407.2
R16 dvss.n1161 dvss.n1148 25407.2
R17 dvss.n786 dvss.n784 25407.2
R18 dvss.n1148 dvss.n784 25407.2
R19 dvss.n1164 dvss.n782 25407.2
R20 dvss.n1164 dvss.n783 25407.2
R21 dvss.n1166 dvss.n782 25407.2
R22 dvss.n1166 dvss.n783 25407.2
R23 dvss.n1277 dvss.n1276 23251
R24 dvss.n1264 dvss.n1259 22647.7
R25 dvss.n896 dvss.n884 21160.1
R26 dvss.n1060 dvss.n884 21160.1
R27 dvss.n896 dvss.n885 21160.1
R28 dvss.n1060 dvss.n885 21160.1
R29 dvss.n1276 dvss.n1275 20409.5
R30 dvss.n1310 dvss.n1309 20031.7
R31 dvss.n1136 dvss.n1135 18221.7
R32 dvss.n1016 dvss.n927 16351
R33 dvss.n1016 dvss.n928 16351
R34 dvss.n968 dvss.n928 16351
R35 dvss.n976 dvss.n790 14459.8
R36 dvss.n1414 dvss.n1413 13403.5
R37 dvss.n1415 dvss.t426 13207.5
R38 dvss.n536 dvss.n48 11399
R39 dvss.n293 dvss.n292 11392.7
R40 dvss.n553 dvss.n552 10626
R41 dvss.n1412 dvss.n25 10590.9
R42 dvss.n1311 dvss.n1310 10051.9
R43 dvss.n463 dvss.n458 9608.16
R44 dvss.n1090 dvss.n838 9322.74
R45 dvss.n1090 dvss.n839 9322.74
R46 dvss.n1102 dvss.n839 9322.74
R47 dvss.n1102 dvss.n838 9322.74
R48 dvss.n464 dvss.n459 9270.59
R49 dvss.n495 dvss.n459 9270.59
R50 dvss.n464 dvss.n460 9270.59
R51 dvss.n495 dvss.n460 9270.59
R52 dvss.n455 dvss.n368 9270.59
R53 dvss.n375 dvss.n368 9270.59
R54 dvss.n455 dvss.n369 9270.59
R55 dvss.n375 dvss.n369 9270.59
R56 dvss.n458 dvss.n457 9139.67
R57 dvss.n1050 dvss.n892 9038.82
R58 dvss.n1050 dvss.n893 9038.82
R59 dvss.n895 dvss.n892 9038.82
R60 dvss.n895 dvss.n893 9038.82
R61 dvss.n754 dvss.n753 9007.72
R62 dvss.n754 dvss.n49 8323.52
R63 dvss.n1066 dvss.n866 8190.47
R64 dvss.n1135 dvss.n790 8011.88
R65 dvss.n1413 dvss.n1412 7594.98
R66 dvss.n1275 dvss.n1260 7497.54
R67 dvss.n1311 dvss.n48 6982.95
R68 dvss.n978 dvss.n788 5937.98
R69 dvss.n878 dvss.n866 5683.2
R70 dvss.n1415 dvss.n1414 5423.26
R71 dvss.n1378 dvss.n29 5288.89
R72 dvss.n936 dvss.n931 5168.35
R73 dvss.n1007 dvss.n936 5168.35
R74 dvss.n1041 dvss.n904 5168.35
R75 dvss.n1029 dvss.n904 5168.35
R76 dvss.n1157 dvss.n1149 5140.55
R77 dvss.n638 dvss 4834.33
R78 dvss.n1137 dvss.n1136 4750.72
R79 dvss.n603 dvss.n602 4692.56
R80 dvss.n966 dvss.n928 4473.2
R81 dvss.n858 dvss.n857 4439.33
R82 dvss.n1297 dvss.n68 4152.6
R83 dvss.n1296 dvss.n68 4152.6
R84 dvss.n880 dvss.n869 4131.21
R85 dvss.n1063 dvss.n869 4131.21
R86 dvss.n880 dvss.n870 4131.21
R87 dvss.n1063 dvss.n870 4131.21
R88 dvss.n639 dvss 4092.31
R89 dvss.n1077 dvss.n1076 4025.74
R90 dvss.n1135 dvss.n1134 4018.37
R91 dvss.n1264 dvss.n1260 3860.74
R92 dvss.n922 dvss.n899 3760.38
R93 dvss.n923 dvss.n922 3760.38
R94 dvss.n1025 dvss.n898 3760.38
R95 dvss.n1025 dvss.n921 3760.38
R96 dvss.n1012 dvss.n1011 3760.38
R97 dvss.n1011 dvss.n933 3760.38
R98 dvss.n967 dvss.n927 3618.97
R99 dvss.n602 dvss.n601 3396.49
R100 dvss.n1087 dvss.n1086 3115.28
R101 dvss.n1087 dvss.n846 3115.28
R102 dvss.n819 dvss.n817 3115.28
R103 dvss.n1124 dvss.n817 3115.28
R104 dvss.n959 dvss.n955 3115.28
R105 dvss.n959 dvss.n957 3115.28
R106 dvss.n847 dvss.n846 3098.81
R107 dvss.n1086 dvss.n847 3098.81
R108 dvss.n1146 dvss.n790 3089.77
R109 dvss.n1307 dvss.n52 3075.76
R110 dvss.n1307 dvss.n51 3075.76
R111 dvss.n1296 dvss.n57 2953.91
R112 dvss.n1297 dvss.n63 2953.91
R113 dvss.n510 dvss.n507 2933.33
R114 dvss.n1146 dvss.n1145 2634.65
R115 dvss.n876 dvss.n854 2575.21
R116 dvss.n876 dvss.n855 2575.21
R117 dvss.n1079 dvss.n855 2575.21
R118 dvss.n1079 dvss.n854 2575.21
R119 dvss.n947 dvss.n806 2575.21
R120 dvss.n1132 dvss.n806 2575.21
R121 dvss.n1132 dvss.n807 2575.21
R122 dvss.n947 dvss.n807 2575.21
R123 dvss.n994 dvss.n942 2575.21
R124 dvss.n999 dvss.n942 2575.21
R125 dvss.n1004 dvss.n938 2575.21
R126 dvss.n1004 dvss.n939 2575.21
R127 dvss.n975 dvss.n789 2476.23
R128 dvss.n976 dvss.n975 2476.23
R129 dvss.n1410 dvss.n1409 2449.56
R130 dvss.n757 dvss.n737 2445.12
R131 dvss.n739 dvss.n737 2445.12
R132 dvss.n765 dvss.n84 2445.12
R133 dvss.n767 dvss.n84 2445.12
R134 dvss.n748 dvss.n740 2445.12
R135 dvss.n748 dvss.n741 2445.12
R136 dvss.n1417 dvss.n1416 2445.12
R137 dvss.n1416 dvss.n22 2445.12
R138 dvss.n978 dvss.n971 2390.79
R139 dvss.n978 dvss.n977 2390.79
R140 dvss.n977 dvss.n974 2390.79
R141 dvss.n974 dvss.n971 2390.79
R142 dvss.n504 dvss.n497 2317.65
R143 dvss.n504 dvss.n501 2317.65
R144 dvss.n1407 dvss.n1379 2317.65
R145 dvss.n1407 dvss.n1380 2317.65
R146 dvss.n1409 dvss.n1378 2284.88
R147 dvss.n1146 dvss.n789 2229.6
R148 dvss.n1121 dvss.n821 2216.26
R149 dvss.n1121 dvss.n818 2216.26
R150 dvss.n539 dvss.n365 2127.34
R151 dvss.n513 dvss.n365 2127.34
R152 dvss.n852 dvss.n850 2064.78
R153 dvss.n1083 dvss.n850 2064.78
R154 dvss.n1083 dvss.n849 2064.78
R155 dvss.n852 dvss.n849 2064.78
R156 dvss.n534 dvss.n514 2016.35
R157 dvss.n534 dvss.n515 2016.35
R158 dvss.n526 dvss.n523 2016.35
R159 dvss.n523 dvss.n522 2016.35
R160 dvss.n649 dvss.n645 2016.35
R161 dvss.n649 dvss.n646 2016.35
R162 dvss.n650 dvss.n645 2016.35
R163 dvss.n650 dvss.n646 2016.35
R164 dvss.n56 dvss.n52 1877.07
R165 dvss.n62 dvss.n51 1877.07
R166 dvss.n421 dvss.n420 1863.9
R167 dvss.n420 dvss.n416 1863.9
R168 dvss.n403 dvss.n366 1863.9
R169 dvss.n412 dvss.n366 1863.9
R170 dvss.n996 dvss.n995 1857.31
R171 dvss.n996 dvss.n943 1857.31
R172 dvss.n550 dvss.n354 1834.26
R173 dvss.n550 dvss.n353 1834.26
R174 dvss.n1280 dvss.n1255 1772.77
R175 dvss.n72 dvss.n69 1735.47
R176 dvss.n72 dvss.n70 1735.47
R177 dvss.n76 dvss.n70 1735.47
R178 dvss.n76 dvss.n69 1735.47
R179 dvss.n1279 dvss.n1256 1653.19
R180 dvss.n1167 dvss.n781 1650.89
R181 dvss.n1160 dvss.n1159 1650.82
R182 dvss.n802 dvss.n798 1603.74
R183 dvss.n1139 dvss.n798 1603.74
R184 dvss.n1144 dvss.n793 1603.74
R185 dvss.n1144 dvss.n792 1603.74
R186 dvss.n1106 dvss.n1105 1603.74
R187 dvss.n1105 dvss.n836 1603.74
R188 dvss.n918 dvss.n910 1603.74
R189 dvss.n918 dvss.n909 1603.74
R190 dvss.n1412 dvss.n1411 1550.2
R191 dvss.n1413 dvss.n27 1539.06
R192 dvss.n1012 dvss.n931 1407.97
R193 dvss.n1013 dvss.n1012 1407.97
R194 dvss.n1013 dvss.n898 1407.97
R195 dvss.n1046 dvss.n898 1407.97
R196 dvss.n1046 dvss.n899 1407.97
R197 dvss.n1041 dvss.n899 1407.97
R198 dvss.n1007 dvss.n933 1407.97
R199 dvss.n933 dvss.n932 1407.97
R200 dvss.n932 dvss.n921 1407.97
R201 dvss.n1033 dvss.n921 1407.97
R202 dvss.n1033 dvss.n923 1407.97
R203 dvss.n1029 dvss.n923 1407.97
R204 dvss.n757 dvss.n95 1344.24
R205 dvss.n739 dvss.n90 1344.24
R206 dvss.n765 dvss.n86 1344.24
R207 dvss.n740 dvss.n86 1344.24
R208 dvss.n767 dvss.n85 1344.24
R209 dvss.n741 dvss.n85 1344.24
R210 dvss.n1424 dvss.n8 1344.24
R211 dvss.n1424 dvss.n20 1344.24
R212 dvss.n1417 dvss.n20 1344.24
R213 dvss.n1426 dvss.n12 1344.24
R214 dvss.n1426 dvss.n19 1344.24
R215 dvss.n22 dvss.n19 1344.24
R216 dvss.n879 dvss.n878 1316.44
R217 dvss.n1273 dvss.n1256 1305.96
R218 dvss.n507 dvss.n506 1303.03
R219 dvss.n920 dvss.n919 1271.1
R220 dvss.n988 dvss.n987 1254.4
R221 dvss.n1061 dvss.n883 1249.02
R222 dvss.n497 dvss.n98 1216.76
R223 dvss.n732 dvss.n98 1216.76
R224 dvss.n732 dvss.n94 1216.76
R225 dvss.n501 dvss.n99 1216.76
R226 dvss.n727 dvss.n99 1216.76
R227 dvss.n727 dvss.n89 1216.76
R228 dvss.n1384 dvss.n1379 1216.76
R229 dvss.n1390 dvss.n1380 1216.76
R230 dvss.n62 dvss.n61 1198.69
R231 dvss.n61 dvss.n56 1198.69
R232 dvss.n65 dvss.n63 1198.69
R233 dvss.n65 dvss.n57 1198.69
R234 dvss.n1168 dvss.n1167 1172.15
R235 dvss.n506 dvss.n496 1141.23
R236 dvss.n372 dvss.n360 1132.83
R237 dvss.n372 dvss.n358 1132.83
R238 dvss.n508 dvss.n361 1132.83
R239 dvss.n508 dvss.n359 1132.83
R240 dvss.n506 dvss.n505 1120.97
R241 dvss.n528 dvss.n519 1100.88
R242 dvss.n528 dvss.n520 1100.88
R243 dvss.n728 dvss.n94 1100.88
R244 dvss.n728 dvss.n89 1100.88
R245 dvss.n498 dvss.n98 1100.88
R246 dvss.n498 dvss.n99 1100.88
R247 dvss.n751 dvss.n95 1100.88
R248 dvss.n751 dvss.n90 1100.88
R249 dvss.n92 dvss.n86 1100.88
R250 dvss.n92 dvss.n85 1100.88
R251 dvss.n16 dvss.n8 1100.88
R252 dvss.n16 dvss.n12 1100.88
R253 dvss.n13 dvss.n7 1100.88
R254 dvss.n13 dvss.n11 1100.88
R255 dvss.n1393 dvss.n1385 1100.88
R256 dvss.n1393 dvss.n1391 1100.88
R257 dvss.n1389 dvss.n1384 1100.88
R258 dvss.n1390 dvss.n1389 1100.88
R259 dvss.n1420 dvss.n20 1100.88
R260 dvss.n1420 dvss.n19 1100.88
R261 dvss.n1160 dvss.n1149 1075.2
R262 dvss.n1272 dvss.n1262 1045.38
R263 dvss.n1038 dvss.n906 1034.77
R264 dvss.n1034 dvss.n920 1033.54
R265 dvss.n1104 dvss.n1103 1032.48
R266 dvss.n404 dvss.n403 994.518
R267 dvss.n430 dvss.n404 994.518
R268 dvss.n430 dvss.n405 994.518
R269 dvss.n416 dvss.n405 994.518
R270 dvss.n412 dvss.n406 994.518
R271 dvss.n428 dvss.n406 994.518
R272 dvss.n428 dvss.n407 994.518
R273 dvss.n421 dvss.n407 994.518
R274 dvss.n545 dvss.n358 994.518
R275 dvss.n545 dvss.n359 994.518
R276 dvss.n513 dvss.n359 994.518
R277 dvss.n543 dvss.n360 994.518
R278 dvss.n543 dvss.n361 994.518
R279 dvss.n539 dvss.n361 994.518
R280 dvss.n1138 dvss.n1137 960.768
R281 dvss.n1159 dvss.n1158 926.37
R282 dvss.n602 dvss.n48 922.37
R283 dvss.n519 dvss.n514 915.471
R284 dvss.n526 dvss.n519 915.471
R285 dvss.n520 dvss.n515 915.471
R286 dvss.n522 dvss.n520 915.471
R287 dvss.n761 dvss.n94 915.471
R288 dvss.n761 dvss.n95 915.471
R289 dvss.n762 dvss.n89 915.471
R290 dvss.n762 dvss.n90 915.471
R291 dvss.n1402 dvss.n1384 915.471
R292 dvss.n1402 dvss.n1385 915.471
R293 dvss.n1396 dvss.n1385 915.471
R294 dvss.n1396 dvss.n7 915.471
R295 dvss.n1431 dvss.n7 915.471
R296 dvss.n1431 dvss.n8 915.471
R297 dvss.n1401 dvss.n1390 915.471
R298 dvss.n1401 dvss.n1391 915.471
R299 dvss.n1397 dvss.n1391 915.471
R300 dvss.n1397 dvss.n11 915.471
R301 dvss.n1430 dvss.n11 915.471
R302 dvss.n1430 dvss.n12 915.471
R303 dvss.n919 dvss.n908 912.745
R304 dvss.n908 dvss.n829 912.745
R305 dvss.n1112 dvss.n829 912.745
R306 dvss.n1112 dvss.n1111 912.745
R307 dvss.n1111 dvss.n831 912.745
R308 dvss.n1104 dvss.n831 912.745
R309 dvss.n1163 dvss.n781 901.063
R310 dvss.n647 dvss.n29 897.29
R311 dvss.n821 dvss.n819 882.553
R312 dvss.n955 dvss.n821 882.553
R313 dvss.n1124 dvss.n818 882.553
R314 dvss.n957 dvss.n818 882.553
R315 dvss.n409 dvss.n406 869.38
R316 dvss.n409 dvss.n404 869.38
R317 dvss.n424 dvss.n407 869.38
R318 dvss.n424 dvss.n405 869.38
R319 dvss.n801 dvss.n800 869.38
R320 dvss.n800 dvss.n797 869.38
R321 dvss.n912 dvss.n911 869.38
R322 dvss.n912 dvss.n827 869.38
R323 dvss.n1110 dvss.n832 869.38
R324 dvss.n1110 dvss.n828 869.38
R325 dvss.n1309 dvss.n50 857.888
R326 dvss.n1309 dvss.n1308 853.793
R327 dvss.n1410 dvss.n25 852.576
R328 dvss.n1103 dvss.n837 844.274
R329 dvss.n1089 dvss.n837 844.274
R330 dvss.n1145 dvss.n791 834.323
R331 dvss.n1302 dvss.n56 833.155
R332 dvss.n1302 dvss.n57 833.155
R333 dvss.n1301 dvss.n62 833.155
R334 dvss.n1301 dvss.n63 833.155
R335 dvss.n799 dvss.n791 829.418
R336 dvss.n1138 dvss.n799 829.418
R337 dvss.n1266 dvss.n1263 818.081
R338 dvss.t256 dvss.t7 793.134
R339 dvss.n640 dvss.n29 768.981
R340 dvss.n906 dvss.n883 762.323
R341 dvss.t253 dvss.t252 759.143
R342 dvss.n1411 dvss.n28 754.202
R343 dvss.t291 dvss.t282 747.812
R344 dvss.t290 dvss.t291 747.812
R345 dvss.n797 dvss.n793 734.362
R346 dvss.n1139 dvss.n797 734.362
R347 dvss.n801 dvss.n792 734.362
R348 dvss.n802 dvss.n801 734.362
R349 dvss.n910 dvss.n827 734.362
R350 dvss.n1113 dvss.n827 734.362
R351 dvss.n1113 dvss.n828 734.362
R352 dvss.n836 dvss.n828 734.362
R353 dvss.n911 dvss.n909 734.362
R354 dvss.n911 dvss.n830 734.362
R355 dvss.n832 dvss.n830 734.362
R356 dvss.n1106 dvss.n832 734.362
R357 dvss.n1313 dvss 719.574
R358 dvss.n995 dvss.n994 717.898
R359 dvss.n995 dvss.n938 717.898
R360 dvss.n999 dvss.n943 717.898
R361 dvss.n943 dvss.n939 717.898
R362 dvss.n1409 dvss.n1408 712.615
R363 dvss.n358 dvss.n354 701.432
R364 dvss.n360 dvss.n353 701.432
R365 dvss.n292 dvss.n158 692.46
R366 dvss.n286 dvss.n285 692.46
R367 dvss.n278 dvss.n178 692.46
R368 dvss.n277 dvss.n276 692.46
R369 dvss.n270 dvss.n269 692.46
R370 dvss.n268 dvss.n192 692.46
R371 dvss.n261 dvss.n260 692.46
R372 dvss.n254 dvss.n253 692.46
R373 dvss.n252 dvss.n222 692.46
R374 dvss.n245 dvss.n244 692.46
R375 dvss.n604 dvss.n115 692.46
R376 dvss.n536 dvss.n535 688.947
R377 dvss.n638 dvss.t255 683.606
R378 dvss.n284 dvss.t309 670.821
R379 dvss.t313 dvss.n221 670.821
R380 dvss.n1005 dvss.n907 640.116
R381 dvss.n1163 dvss.n780 639.551
R382 dvss.n1123 dvss.n805 634.548
R383 dvss.n958 dvss.n820 634.548
R384 dvss.n262 dvss.t374 627.542
R385 dvss.t317 dvss.n603 627.542
R386 dvss.t430 dvss.t263 626.923
R387 dvss.n1123 dvss.n1122 622.928
R388 dvss.n1122 dvss.n820 622.928
R389 dvss.n987 dvss.n986 620.308
R390 dvss.n1377 dvss.n1376 611.778
R391 dvss.n1315 dvss.n1314 611.778
R392 dvss.n641 dvss.n640 611.778
R393 dvss.n709 dvss.n47 611.778
R394 dvss.n537 dvss.n536 599.069
R395 dvss.n376 dvss.n371 594.447
R396 dvss.n494 dvss.n461 594.447
R397 dvss.n291 dvss.n290 585
R398 dvss.n292 dvss.n291 585
R399 dvss.n289 dvss.n159 585
R400 dvss.n159 dvss.n158 585
R401 dvss.n288 dvss.n287 585
R402 dvss.n287 dvss.n286 585
R403 dvss.n166 dvss.n165 585
R404 dvss.n285 dvss.n166 585
R405 dvss.n283 dvss.n282 585
R406 dvss.n284 dvss.n283 585
R407 dvss.n281 dvss.n167 585
R408 dvss.n178 dvss.n167 585
R409 dvss.n280 dvss.n279 585
R410 dvss.n279 dvss.n278 585
R411 dvss.n177 dvss.n176 585
R412 dvss.n277 dvss.n177 585
R413 dvss.n275 dvss.n274 585
R414 dvss.n276 dvss.n275 585
R415 dvss.n273 dvss.n179 585
R416 dvss.n191 dvss.n179 585
R417 dvss.n272 dvss.n271 585
R418 dvss.n271 dvss.n270 585
R419 dvss.n190 dvss.n189 585
R420 dvss.n269 dvss.n190 585
R421 dvss.n267 dvss.n266 585
R422 dvss.n268 dvss.n267 585
R423 dvss.n265 dvss.n193 585
R424 dvss.n193 dvss.n192 585
R425 dvss.n264 dvss.n263 585
R426 dvss.n263 dvss.n262 585
R427 dvss.n204 dvss.n203 585
R428 dvss.n261 dvss.n204 585
R429 dvss.n259 dvss.n258 585
R430 dvss.n260 dvss.n259 585
R431 dvss.n257 dvss.n205 585
R432 dvss.n221 dvss.n205 585
R433 dvss.n256 dvss.n255 585
R434 dvss.n255 dvss.n254 585
R435 dvss.n220 dvss.n219 585
R436 dvss.n253 dvss.n220 585
R437 dvss.n251 dvss.n250 585
R438 dvss.n252 dvss.n251 585
R439 dvss.n249 dvss.n223 585
R440 dvss.n223 dvss.n222 585
R441 dvss.n248 dvss.n247 585
R442 dvss.n247 dvss.n246 585
R443 dvss.n234 dvss.n233 585
R444 dvss.n245 dvss.n234 585
R445 dvss.n243 dvss.n242 585
R446 dvss.n244 dvss.n243 585
R447 dvss.n113 dvss.n111 585
R448 dvss.n115 dvss.n113 585
R449 dvss.n606 dvss.n605 585
R450 dvss.n605 dvss.n604 585
R451 dvss.n114 dvss.n112 585
R452 dvss.n603 dvss.n114 585
R453 dvss.n295 dvss.n294 585
R454 dvss.n294 dvss.n293 585
R455 dvss.n301 dvss.n300 585
R456 dvss.n302 dvss.n301 585
R457 dvss.n157 dvss.n156 585
R458 dvss.n303 dvss.n157 585
R459 dvss.n307 dvss.n306 585
R460 dvss.n306 dvss.n305 585
R461 dvss.n152 dvss.n151 585
R462 dvss.n304 dvss.n151 585
R463 dvss.n315 dvss.n314 585
R464 dvss.n315 dvss.n150 585
R465 dvss.n316 dvss.n148 585
R466 dvss.n317 dvss.n316 585
R467 dvss.n323 dvss.n149 585
R468 dvss.n318 dvss.n149 585
R469 dvss.n322 dvss.n321 585
R470 dvss.n321 dvss.n320 585
R471 dvss.n144 dvss.n143 585
R472 dvss.n319 dvss.n143 585
R473 dvss.n336 dvss.n335 585
R474 dvss.n337 dvss.n336 585
R475 dvss.n142 dvss.n141 585
R476 dvss.n338 dvss.n142 585
R477 dvss.n342 dvss.n341 585
R478 dvss.n341 dvss.n340 585
R479 dvss.n137 dvss.n136 585
R480 dvss.n339 dvss.n136 585
R481 dvss.n350 dvss.n349 585
R482 dvss.n351 dvss.n350 585
R483 dvss.n135 dvss.n134 585
R484 dvss.n352 dvss.n135 585
R485 dvss.n557 dvss.n556 585
R486 dvss.n556 dvss.n555 585
R487 dvss.n130 dvss.n129 585
R488 dvss.n554 dvss.n129 585
R489 dvss.n565 dvss.n564 585
R490 dvss.n565 dvss.n128 585
R491 dvss.n566 dvss.n126 585
R492 dvss.n567 dvss.n566 585
R493 dvss.n573 dvss.n127 585
R494 dvss.n568 dvss.n127 585
R495 dvss.n572 dvss.n571 585
R496 dvss.n571 dvss.n570 585
R497 dvss.n122 dvss.n121 585
R498 dvss.n569 dvss.n121 585
R499 dvss.n586 dvss.n585 585
R500 dvss.n587 dvss.n586 585
R501 dvss.n120 dvss.n119 585
R502 dvss.n588 dvss.n120 585
R503 dvss.n592 dvss.n591 585
R504 dvss.n591 dvss.n590 585
R505 dvss.n117 dvss.n116 585
R506 dvss.n589 dvss.n116 585
R507 dvss.n600 dvss.n599 585
R508 dvss.n601 dvss.n600 585
R509 dvss.t134 dvss.n191 584.263
R510 dvss.n246 dvss.t25 584.263
R511 dvss.n1088 dvss.n845 580.571
R512 dvss.n1076 dvss.n857 576
R513 dvss.n1036 dvss.n845 569.938
R514 dvss.n1082 dvss.n851 559.304
R515 dvss.n1082 dvss.n1081 559.304
R516 dvss.t282 dvss.n47 555.193
R517 dvss.n466 dvss.n461 554.4
R518 dvss.n453 dvss.n371 554.201
R519 dvss.t180 dvss.n1377 543.211
R520 dvss.n1035 dvss.n1034 542.292
R521 dvss.n191 dvss.t94 540.985
R522 dvss.n246 dvss.t16 540.985
R523 dvss.n291 dvss.n159 539.294
R524 dvss.n287 dvss.n159 539.294
R525 dvss.n287 dvss.n166 539.294
R526 dvss.n283 dvss.n166 539.294
R527 dvss.n283 dvss.n167 539.294
R528 dvss.n279 dvss.n167 539.294
R529 dvss.n279 dvss.n177 539.294
R530 dvss.n275 dvss.n177 539.294
R531 dvss.n275 dvss.n179 539.294
R532 dvss.n271 dvss.n179 539.294
R533 dvss.n271 dvss.n190 539.294
R534 dvss.n267 dvss.n190 539.294
R535 dvss.n267 dvss.n193 539.294
R536 dvss.n263 dvss.n193 539.294
R537 dvss.n263 dvss.n204 539.294
R538 dvss.n259 dvss.n204 539.294
R539 dvss.n259 dvss.n205 539.294
R540 dvss.n255 dvss.n205 539.294
R541 dvss.n255 dvss.n220 539.294
R542 dvss.n251 dvss.n220 539.294
R543 dvss.n251 dvss.n223 539.294
R544 dvss.n247 dvss.n223 539.294
R545 dvss.n247 dvss.n234 539.294
R546 dvss.n243 dvss.n234 539.294
R547 dvss.n243 dvss.n113 539.294
R548 dvss.n605 dvss.n113 539.294
R549 dvss.n605 dvss.n114 539.294
R550 dvss.n301 dvss.n294 539.294
R551 dvss.n301 dvss.n157 539.294
R552 dvss.n306 dvss.n157 539.294
R553 dvss.n306 dvss.n151 539.294
R554 dvss.n315 dvss.n151 539.294
R555 dvss.n316 dvss.n315 539.294
R556 dvss.n316 dvss.n149 539.294
R557 dvss.n321 dvss.n149 539.294
R558 dvss.n321 dvss.n143 539.294
R559 dvss.n336 dvss.n143 539.294
R560 dvss.n336 dvss.n142 539.294
R561 dvss.n341 dvss.n142 539.294
R562 dvss.n341 dvss.n136 539.294
R563 dvss.n350 dvss.n136 539.294
R564 dvss.n350 dvss.n135 539.294
R565 dvss.n556 dvss.n135 539.294
R566 dvss.n556 dvss.n129 539.294
R567 dvss.n565 dvss.n129 539.294
R568 dvss.n566 dvss.n565 539.294
R569 dvss.n566 dvss.n127 539.294
R570 dvss.n571 dvss.n127 539.294
R571 dvss.n571 dvss.n121 539.294
R572 dvss.n586 dvss.n121 539.294
R573 dvss.n586 dvss.n120 539.294
R574 dvss.n591 dvss.n120 539.294
R575 dvss.n591 dvss.n116 539.294
R576 dvss.n600 dvss.n116 539.294
R577 dvss.n77 dvss.t237 538.484
R578 dvss.t237 dvss.n27 538.484
R579 dvss.n881 dvss.n871 538.038
R580 dvss.n1100 dvss.n841 532.726
R581 dvss.t377 dvss.n59 518.009
R582 dvss.t377 dvss.n60 518.009
R583 dvss.n804 dvss.n803 506.709
R584 dvss.n998 dvss.n944 498.207
R585 dvss.t64 dvss.n158 497.705
R586 dvss.n262 dvss.t136 497.705
R587 dvss.n1308 dvss.t422 497.534
R588 dvss.n59 dvss.t424 497.534
R589 dvss.t208 dvss.n60 497.534
R590 dvss.t183 dvss.n78 497.534
R591 dvss.n1035 dvss.n907 491.252
R592 dvss.n1298 dvss.n67 479.248
R593 dvss.n958 dvss.n944 474.168
R594 dvss.t250 dvss.n647 471.003
R595 dvss.t250 dvss.n28 471.003
R596 dvss.n1080 dvss.n853 463.606
R597 dvss.n871 dvss.n853 463.606
R598 dvss.n998 dvss.n997 463.606
R599 dvss.n997 dvss.n937 463.606
R600 dvss.t222 dvss.n284 454.426
R601 dvss.n221 dvss.t68 454.426
R602 dvss.n463 dvss.t297 447.74
R603 dvss.n496 dvss.t234 447.74
R604 dvss.t379 dvss.t422 446.348
R605 dvss.t424 dvss.t88 446.348
R606 dvss.t171 dvss.t208 446.348
R607 dvss.t224 dvss.t171 446.348
R608 dvss.t228 dvss.t224 446.348
R609 dvss.t228 dvss.t115 446.348
R610 dvss.t115 dvss.t19 446.348
R611 dvss.t19 dvss.t183 446.348
R612 dvss.n1134 dvss.n1133 443.952
R613 dvss.n1158 dvss.n1157 443.057
R614 dvss.n457 dvss.t30 442.741
R615 dvss.n1089 dvss.n1088 442.339
R616 dvss.n878 dvss.n857 440.32
R617 dvss.n509 dvss.t10 436.089
R618 dvss.t50 dvss.n537 436.089
R619 dvss dvss.t180 434.568
R620 dvss.t155 dvss.t143 430.558
R621 dvss.t147 dvss.t149 430.558
R622 dvss.n1268 dvss.n1267 426.846
R623 dvss.t141 dvss 426.781
R624 dvss.n1378 dvss 423.252
R625 dvss.t7 dvss.t253 415.452
R626 dvss.n278 dvss.t295 411.149
R627 dvss.n253 dvss.t66 411.149
R628 dvss.t368 dvss 405.144
R629 dvss.t260 dvss.n639 404.12
R630 dvss.n1133 dvss.n805 402.113
R631 dvss.n1085 dvss.n841 401.372
R632 dvss.n1006 dvss.n1005 393.428
R633 dvss.n570 dvss.n568 390.029
R634 dvss.n588 dvss.n587 390.029
R635 dvss.n590 dvss.n589 390.029
R636 dvss.n870 dvss.n866 387.457
R637 dvss dvss.t413 385.236
R638 dvss.t73 dvss.t258 385.236
R639 dvss.t398 dvss.n10 384.057
R640 dvss.n1419 dvss.t401 384.057
R641 dvss.n1419 dvss.t428 384.057
R642 dvss.n1039 dvss.n1038 381.606
R643 dvss.n1101 dvss.n1100 381.137
R644 dvss.t252 dvss.t264 377.683
R645 dvss.t145 dvss.t153 377.683
R646 dvss dvss.t284 373.906
R647 dvss.n302 dvss.n293 371.505
R648 dvss.n305 dvss.n303 371.505
R649 dvss.n317 dvss.n150 371.505
R650 dvss.n320 dvss.n318 371.505
R651 dvss.n338 dvss.n337 371.505
R652 dvss.n340 dvss.n339 371.505
R653 dvss.n555 dvss.n352 371.505
R654 dvss.n567 dvss.n128 371.505
R655 dvss.n882 dvss.n881 367.908
R656 dvss.n1062 dvss.n882 367.908
R657 dvss.t86 dvss.n268 367.87
R658 dvss.t23 dvss.n115 367.87
R659 dvss.n1345 dvss.t114 367.125
R660 dvss.n1414 dvss.n26 364.601
R661 dvss.n304 dvss.t372 359.894
R662 dvss.t5 dvss.t368 359.877
R663 dvss.n1408 dvss.t320 359.637
R664 dvss.n1387 dvss.t322 359.637
R665 dvss.t284 dvss.t288 358.798
R666 dvss.n1306 dvss.n53 356.142
R667 dvss.n601 dvss.t54 353.464
R668 dvss.t2 dvss.n1387 350.757
R669 dvss.t2 dvss.n1388 350.757
R670 dvss.t394 dvss.n1388 350.757
R671 dvss.t394 dvss.n9 350.757
R672 dvss.t44 dvss.n9 350.757
R673 dvss.t44 dvss.n10 350.757
R674 dvss.n1299 dvss.n1298 337.695
R675 dvss.n351 dvss.t293 336.675
R676 dvss.n753 dvss.n752 335.473
R677 dvss.n505 dvss.t370 331.382
R678 dvss.t109 dvss.n499 331.382
R679 dvss.n499 dvss.t77 331.382
R680 dvss.n569 dvss.t70 329.087
R681 dvss.t143 dvss.t141 328.584
R682 dvss.n750 dvss.n749 325.548
R683 dvss.n1081 dvss.n1080 325.375
R684 dvss.t149 dvss.t155 324.808
R685 dvss.t153 dvss.t147 324.808
R686 dvss.t151 dvss.t145 324.808
R687 dvss.t286 dvss.t151 324.808
R688 dvss.t288 dvss.t286 324.808
R689 dvss.n269 dvss.t86 324.591
R690 dvss.n244 dvss.t23 324.591
R691 dvss.t60 dvss.t111 316.837
R692 dvss.t203 dvss.n93 315.017
R693 dvss.n1085 dvss.n1084 313.601
R694 dvss.n319 dvss.t92 313.457
R695 dvss.n730 dvss.n729 310.925
R696 dvss dvss.t175 307.82
R697 dvss.n535 dvss.t48 304.913
R698 dvss.n527 dvss.t48 304.913
R699 dvss.n527 dvss.t388 304.913
R700 dvss.t388 dvss.n521 304.913
R701 dvss.n951 dvss.n950 304.849
R702 dvss.t130 dvss.n569 304.709
R703 dvss.t52 dvss.n510 299.2
R704 dvss.t18 dvss.t260 294.592
R705 dvss.t264 dvss.t18 294.592
R706 dvss.t413 dvss.t256 294.592
R707 dvss.t255 dvss.t73 294.592
R708 dvss.n1023 dvss.n895 292.5
R709 dvss.n1049 dvss.n895 292.5
R710 dvss.n1051 dvss.n1050 292.5
R711 dvss.n1050 dvss.n1049 292.5
R712 dvss.n1430 dvss.n1429 292.5
R713 dvss.t44 dvss.n1430 292.5
R714 dvss.n1398 dvss.n1397 292.5
R715 dvss.n1397 dvss.t394 292.5
R716 dvss.n1401 dvss.n1400 292.5
R717 dvss.t2 dvss.n1401 292.5
R718 dvss.n1403 dvss.n1402 292.5
R719 dvss.n1402 dvss.t2 292.5
R720 dvss.n1396 dvss.n1395 292.5
R721 dvss.t394 dvss.n1396 292.5
R722 dvss.n1432 dvss.n1431 292.5
R723 dvss.n1431 dvss.t44 292.5
R724 dvss.n651 dvss.n650 292.5
R725 dvss.n650 dvss.t250 292.5
R726 dvss.n649 dvss.n648 292.5
R727 dvss.t250 dvss.n649 292.5
R728 dvss.n522 dvss.n517 292.5
R729 dvss.t388 dvss.n522 292.5
R730 dvss.n532 dvss.n515 292.5
R731 dvss.n515 dvss.t48 292.5
R732 dvss.n516 dvss.n514 292.5
R733 dvss.n514 dvss.t48 292.5
R734 dvss.n526 dvss.n525 292.5
R735 dvss.t388 dvss.n526 292.5
R736 dvss.n763 dvss.n762 292.5
R737 dvss.n762 dvss.t203 292.5
R738 dvss.n761 dvss.n760 292.5
R739 dvss.t203 dvss.n761 292.5
R740 dvss.t138 dvss.n319 290.238
R741 dvss.n78 dvss.n77 286.646
R742 dvss.n553 dvss.t0 286.368
R743 dvss.t295 dvss.n277 281.312
R744 dvss.t66 dvss.n252 281.312
R745 dvss.n1368 dvss.t481 280.997
R746 dvss.n1053 dvss.n886 274.389
R747 dvss.n1354 dvss.t176 274.164
R748 dvss.t258 dvss.t290 271.932
R749 dvss.n1411 dvss.n1410 271.274
R750 dvss.n374 dvss.n373 268.997
R751 dvss.t21 dvss.n302 267.019
R752 dvss.t14 dvss.n351 267.019
R753 dvss.t297 dvss.t96 265.327
R754 dvss.t96 dvss.t164 265.327
R755 dvss.t164 dvss.t230 265.327
R756 dvss.t230 dvss.t405 265.327
R757 dvss.t405 dvss.t98 265.327
R758 dvss.t98 dvss.t232 265.327
R759 dvss.t232 dvss.t301 265.327
R760 dvss.t301 dvss.t307 265.327
R761 dvss.t307 dvss.t384 265.327
R762 dvss.t384 dvss.t433 265.327
R763 dvss.t433 dvss.t403 265.327
R764 dvss.t403 dvss.t299 265.327
R765 dvss.t299 dvss.t119 265.327
R766 dvss.t119 dvss.t162 265.327
R767 dvss.t162 dvss.t303 265.327
R768 dvss.t303 dvss.t267 265.327
R769 dvss.t267 dvss.t56 265.327
R770 dvss.t56 dvss.t277 265.327
R771 dvss.t277 dvss.t269 265.327
R772 dvss.t269 dvss.t273 265.327
R773 dvss.t273 dvss.t58 265.327
R774 dvss.t58 dvss.t271 265.327
R775 dvss.t271 dvss.t275 265.327
R776 dvss.t275 dvss.t336 265.327
R777 dvss.t336 dvss.t334 265.327
R778 dvss.t334 dvss.t234 265.327
R779 dvss.n1136 dvss.n803 262.652
R780 dvss.t175 dvss.t37 258.026
R781 dvss.n676 dvss.t257 255.72
R782 dvss.n454 dvss.n370 252.941
R783 dvss.n465 dvss.n462 252.941
R784 dvss.n1375 dvss.t181 251.179
R785 dvss.n540 dvss.n364 247.719
R786 dvss.n703 dvss.t292 246.01
R787 dvss.n1010 dvss.n934 244.329
R788 dvss.n1010 dvss.n1009 244.329
R789 dvss.n1043 dvss.n902 244.329
R790 dvss.n1031 dvss.n902 244.329
R791 dvss.n1026 dvss.n1024 244.329
R792 dvss.n1027 dvss.n1026 244.329
R793 dvss.t132 dvss.n304 243.799
R794 dvss.t218 dvss.n554 243.799
R795 dvss.n966 dvss.n965 238.726
R796 dvss.n285 dvss.t222 238.034
R797 dvss.n260 dvss.t68 238.034
R798 dvss.t412 dvss 237.655
R799 dvss.n384 dvss.t80 236.52
R800 dvss.n473 dvss.t298 236.52
R801 dvss.n716 dvss.t371 236.333
R802 dvss.n719 dvss.t206 236.3
R803 dvss.n721 dvss.t78 236.243
R804 dvss.n721 dvss.t110 236.212
R805 dvss.t113 dvss.t166 235.535
R806 dvss.n717 dvss.t351 231.785
R807 dvss.n106 dvss.t389 231.564
R808 dvss.n2 dvss.t395 231.562
R809 dvss.n3 dvss.t45 231.562
R810 dvss.n1 dvss.t3 231.56
R811 dvss.n107 dvss.t49 231.554
R812 dvss.n771 dvss.t408 231.512
R813 dvss.n642 dvss.t251 231.501
R814 dvss.n772 dvss.t202 231.401
R815 dvss.n718 dvss.t204 231.357
R816 dvss.n717 dvss.t366 231.351
R817 dvss.t420 dvss.t419 230.934
R818 dvss.t280 dvss.t5 230.864
R819 dvss.n1335 dvss.n1334 230.579
R820 dvss.n961 dvss.n953 227.097
R821 dvss.n1368 dvss.t182 223.571
R822 dvss.n58 dvss.t379 223.174
R823 dvss.t88 dvss.n58 223.174
R824 dvss.t265 dvss.n317 220.581
R825 dvss.n991 dvss.n940 216.847
R826 dvss.n965 dvss.n964 215.651
R827 dvss.n964 dvss.n929 215.651
R828 dvss.n1040 dvss.n905 215.651
R829 dvss.n1040 dvss.n1039 215.651
R830 dvss.n1348 dvss.n1347 215.293
R831 dvss.n64 dvss.n53 214.589
R832 dvss.n549 dvss.n355 214.213
R833 dvss.t216 dvss.n567 213.03
R834 dvss.n624 dvss.n623 212.733
R835 dvss.n1059 dvss.n1058 211.93
R836 dvss.n635 dvss.n634 211.183
R837 dvss.n657 dvss.n637 211.183
R838 dvss.n1295 dvss.n67 210.745
R839 dvss.n1001 dvss.n940 210.447
R840 dvss.n755 dvss.n750 209.524
R841 dvss.n669 dvss.n628 209.243
R842 dvss.n631 dvss.n630 209.243
R843 dvss.n663 dvss.n633 209.243
R844 dvss.n617 dvss.n616 208.856
R845 dvss.n968 dvss.n967 208.383
R846 dvss.n590 dvss.t128 207.202
R847 dvss.n1310 dvss.n49 206.857
R848 dvss.n43 dvss.n42 206.528
R849 dvss.n1037 dvss.n851 206.284
R850 dvss.n690 dvss.n689 205.282
R851 dvss.t340 dvss.t32 205.274
R852 dvss.t392 dvss.t199 204.95
R853 dvss.t390 dvss.t438 204.95
R854 dvss.t214 dvss.t390 204.95
R855 dvss.t386 dvss.t212 204.95
R856 dvss.n73 dvss.n71 202.918
R857 dvss.n74 dvss.n73 202.918
R858 dvss.n75 dvss.n74 202.918
R859 dvss.n75 dvss.n71 202.918
R860 dvss.t220 dvss.t392 202.796
R861 dvss.t102 dvss.t79 202.397
R862 dvss.t42 dvss.t100 202.397
R863 dvss.t100 dvss.t189 202.397
R864 dvss.t191 dvss.t185 202.397
R865 dvss.t381 dvss.t191 202.397
R866 dvss.t104 dvss.t187 202.397
R867 dvss.t46 dvss.t168 202.397
R868 dvss.t40 dvss.t240 202.397
R869 dvss.t240 dvss.t226 202.397
R870 dvss.t90 dvss.t220 202.397
R871 dvss.n340 dvss.t311 197.362
R872 dvss.n1 dvss.n0 197.084
R873 dvss.n1153 dvss.n1150 196.851
R874 dvss.n1152 dvss.n1151 196.849
R875 dvss.n444 dvss.n443 196.792
R876 dvss.n445 dvss.n395 196.763
R877 dvss.n446 dvss.n394 196.763
R878 dvss.n447 dvss.n393 196.763
R879 dvss.n448 dvss.n392 196.763
R880 dvss.n449 dvss.n391 196.763
R881 dvss.n450 dvss.n390 196.763
R882 dvss.n389 dvss.n378 196.763
R883 dvss.n388 dvss.n379 196.763
R884 dvss.n387 dvss.n380 196.763
R885 dvss.n386 dvss.n381 196.763
R886 dvss.n385 dvss.n382 196.763
R887 dvss.n384 dvss.n383 196.763
R888 dvss.n473 dvss.n472 196.763
R889 dvss.n474 dvss.n471 196.763
R890 dvss.n475 dvss.n470 196.763
R891 dvss.n476 dvss.n469 196.763
R892 dvss.n477 dvss.n468 196.763
R893 dvss.n478 dvss.n467 196.763
R894 dvss.n490 dvss.n479 196.763
R895 dvss.n489 dvss.n480 196.763
R896 dvss.n488 dvss.n481 196.763
R897 dvss.n487 dvss.n482 196.763
R898 dvss.n486 dvss.n483 196.763
R899 dvss.n485 dvss.n484 196.763
R900 dvss.n103 dvss.n102 196.763
R901 dvss.n882 dvss.n870 195
R902 dvss.n874 dvss.n869 195
R903 dvss.n882 dvss.n869 195
R904 dvss.n286 dvss.t64 194.755
R905 dvss.t136 dvss.n261 194.755
R906 dvss.t168 dvss.t243 193.964
R907 dvss.t199 dvss.n551 192.141
R908 dvss.n1107 dvss.n834 187.859
R909 dvss.n917 dvss.n915 187.859
R910 dvss.n423 dvss.t104 187.638
R911 dvss.n1084 dvss.n848 186.058
R912 dvss.t128 dvss.n588 182.826
R913 dvss.n1306 dvss.n1305 181.679
R914 dvss.n640 dvss 181.288
R915 dvss.n949 dvss.n948 177.589
R916 dvss.t37 dvss.t280 176.543
R917 dvss.t311 dvss.n338 174.143
R918 dvss.t212 dvss.t158 172.927
R919 dvss.n708 dvss.t283 171.77
R920 dvss.n1313 dvss.t113 168.239
R921 dvss.t75 dvss.n367 166.555
R922 dvss.n429 dvss.t107 166.555
R923 dvss.n1314 dvss.t160 165.113
R924 dvss.n835 dvss.n834 165.014
R925 dvss.n917 dvss.n916 165.014
R926 dvss.n1047 dvss.n897 164.179
R927 dvss.n926 dvss.n889 161.438
R928 dvss.n24 dvss.n23 159.054
R929 dvss.n758 dvss.n736 159.01
R930 dvss.n568 dvss.t216 158.45
R931 dvss.n408 dvss.t102 158.123
R932 dvss.n422 dvss.t210 158.123
R933 dvss.n30 dvss.t369 156.095
R934 dvss.n374 dvss.t12 155.829
R935 dvss.n671 dvss.t142 154.727
R936 dvss.n544 dvss.t12 154.489
R937 dvss.n544 dvss.t10 154.489
R938 dvss.n538 dvss.t52 154.489
R939 dvss.n538 dvss.t50 154.489
R940 dvss.t121 dvss.t305 151.798
R941 dvss.t112 dvss.t61 151.725
R942 dvss.n276 dvss.t94 151.476
R943 dvss.t16 dvss.n222 151.476
R944 dvss.n318 dvss.t265 150.923
R945 dvss.n1406 dvss.n1381 150.399
R946 dvss.n503 dvss.n502 150.398
R947 dvss.n1312 dvss 149.173
R948 dvss.n355 dvss.n353 146.25
R949 dvss.t158 dvss.n353 146.25
R950 dvss.n548 dvss.n354 146.25
R951 dvss.t158 dvss.n354 146.25
R952 dvss.n376 dvss.n375 146.25
R953 dvss.n375 dvss.n374 146.25
R954 dvss.n1107 dvss.n1106 146.25
R955 dvss.n1106 dvss.n831 146.25
R956 dvss.n833 dvss.n830 146.25
R957 dvss.n1112 dvss.n830 146.25
R958 dvss.n915 dvss.n909 146.25
R959 dvss.n909 dvss.n908 146.25
R960 dvss.n836 dvss.n835 146.25
R961 dvss.n836 dvss.n831 146.25
R962 dvss.n1114 dvss.n1113 146.25
R963 dvss.n1113 dvss.n1112 146.25
R964 dvss.n916 dvss.n910 146.25
R965 dvss.n910 dvss.n908 146.25
R966 dvss.n872 dvss.n854 146.25
R967 dvss.n854 dvss.n853 146.25
R968 dvss.n865 dvss.n855 146.25
R969 dvss.n855 dvss.n853 146.25
R970 dvss.n949 dvss.n806 146.25
R971 dvss.n806 dvss.n804 146.25
R972 dvss.n994 dvss.n993 146.25
R973 dvss.n998 dvss.n994 146.25
R974 dvss.n990 dvss.n938 146.25
R975 dvss.n938 dvss.n937 146.25
R976 dvss.n945 dvss.n807 146.25
R977 dvss.n807 dvss.n804 146.25
R978 dvss.n1002 dvss.n939 146.25
R979 dvss.n939 dvss.n937 146.25
R980 dvss.n1000 dvss.n999 146.25
R981 dvss.n999 dvss.n998 146.25
R982 dvss.n809 dvss.n802 146.25
R983 dvss.n1138 dvss.n802 146.25
R984 dvss.n794 dvss.n792 146.25
R985 dvss.n792 dvss.n791 146.25
R986 dvss.n1140 dvss.n1139 146.25
R987 dvss.n1139 dvss.n1138 146.25
R988 dvss.n1142 dvss.n793 146.25
R989 dvss.n793 dvss.n791 146.25
R990 dvss.n1416 dvss.n24 146.25
R991 dvss.n1416 dvss.n1415 146.25
R992 dvss.n1389 dvss.n1382 146.25
R993 dvss.n1389 dvss.n1387 146.25
R994 dvss.n1394 dvss.n1393 146.25
R995 dvss.n1393 dvss.n1388 146.25
R996 dvss.n14 dvss.n13 146.25
R997 dvss.n13 dvss.n9 146.25
R998 dvss.n17 dvss.n16 146.25
R999 dvss.n16 dvss.n10 146.25
R1000 dvss.n1421 dvss.n1420 146.25
R1001 dvss.n1420 dvss.n1419 146.25
R1002 dvss.n1381 dvss.n1380 146.25
R1003 dvss.n1386 dvss.n1380 146.25
R1004 dvss.n1407 dvss.n1406 146.25
R1005 dvss.n1408 dvss.n1407 146.25
R1006 dvss.n1405 dvss.n1379 146.25
R1007 dvss.n1386 dvss.n1379 146.25
R1008 dvss.n646 dvss.n644 146.25
R1009 dvss.n646 dvss.n28 146.25
R1010 dvss.n645 dvss.n643 146.25
R1011 dvss.n647 dvss.n645 146.25
R1012 dvss.n748 dvss.n747 146.25
R1013 dvss.n749 dvss.n748 146.25
R1014 dvss.n737 dvss.n736 146.25
R1015 dvss.n737 dvss.n50 146.25
R1016 dvss.n529 dvss.n528 146.25
R1017 dvss.n528 dvss.n527 146.25
R1018 dvss.n524 dvss.n523 146.25
R1019 dvss.n523 dvss.n521 146.25
R1020 dvss.n534 dvss.n533 146.25
R1021 dvss.n535 dvss.n534 146.25
R1022 dvss.n92 dvss.n91 146.25
R1023 dvss.n93 dvss.n92 146.25
R1024 dvss.n84 dvss.n82 146.25
R1025 dvss.n730 dvss.n84 146.25
R1026 dvss.n498 dvss.n100 146.25
R1027 dvss.n499 dvss.n498 146.25
R1028 dvss.n728 dvss.n96 146.25
R1029 dvss.n729 dvss.n728 146.25
R1030 dvss.n751 dvss.n735 146.25
R1031 dvss.n752 dvss.n751 146.25
R1032 dvss.n727 dvss.n726 146.25
R1033 dvss.n731 dvss.n727 146.25
R1034 dvss.n501 dvss.n101 146.25
R1035 dvss.n501 dvss.n500 146.25
R1036 dvss.n504 dvss.n503 146.25
R1037 dvss.n505 dvss.n504 146.25
R1038 dvss.n502 dvss.n497 146.25
R1039 dvss.n500 dvss.n497 146.25
R1040 dvss.n733 dvss.n732 146.25
R1041 dvss.n732 dvss.n731 146.25
R1042 dvss.n495 dvss.n494 146.25
R1043 dvss.n496 dvss.n495 146.25
R1044 dvss.n465 dvss.n464 146.25
R1045 dvss.n464 dvss.n463 146.25
R1046 dvss.n455 dvss.n454 146.25
R1047 dvss.n456 dvss.n455 146.25
R1048 dvss.n512 dvss.n364 145.726
R1049 dvss.t245 dvss.t239 144.476
R1050 dvss.t157 dvss.t238 144.476
R1051 dvss.t124 dvss.t140 144.476
R1052 dvss.t9 dvss.t242 144.476
R1053 dvss.t342 dvss.t179 144.476
R1054 dvss.t367 dvss.t72 144.476
R1055 dvss.t29 dvss.t34 144.476
R1056 dvss.t106 dvss.t27 144.476
R1057 dvss.t414 dvss.t38 144.476
R1058 dvss.t62 dvss.t432 144.476
R1059 dvss.t400 dvss.t118 144.476
R1060 dvss.t174 dvss.t437 144.476
R1061 dvss.t279 dvss.t178 144.476
R1062 dvss.t339 dvss.t177 144.476
R1063 dvss.t397 dvss.t85 144.476
R1064 dvss.t315 dvss.t249 144.476
R1065 dvss.t316 dvss.t262 144.476
R1066 dvss.t123 dvss.t247 144.476
R1067 dvss.t409 dvss.t28 144.476
R1068 dvss.t173 dvss.t383 144.476
R1069 dvss.t4 dvss.t436 144.476
R1070 dvss.t117 dvss.t435 144.476
R1071 dvss.n1299 dvss.n66 141.554
R1072 dvss.n64 dvss.n54 141.554
R1073 dvss.n549 dvss.n548 140.059
R1074 dvss.n510 dvss.n509 136.889
R1075 dvss.n1015 dvss.n929 136.668
R1076 dvss.n362 dvss.n356 134.024
R1077 dvss.n541 dvss.n363 134.024
R1078 dvss.n952 dvss.n951 133.369
R1079 dvss.n1095 dvss.n840 131.964
R1080 dvss.n1049 dvss.n1048 131.344
R1081 dvss.n1334 dvss.t341 131.141
R1082 dvss.n533 dvss.n516 131.012
R1083 dvss.n525 dvss.n524 131.012
R1084 dvss.n66 dvss.n55 131.012
R1085 dvss.n1304 dvss.n54 131.012
R1086 dvss.n648 dvss.n643 131.012
R1087 dvss.n648 dvss.n644 131.012
R1088 dvss.n1425 dvss.t398 130.98
R1089 dvss.n1425 dvss.t401 130.98
R1090 dvss.t428 dvss.n1418 130.98
R1091 dvss.n1418 dvss.t426 130.98
R1092 dvss.n1143 dvss.n794 130.087
R1093 dvss.n419 dvss.t40 128.607
R1094 dvss.n46 dvss.n45 128.178
R1095 dvss.n305 dvss.t132 127.704
R1096 dvss.n555 dvss.t218 127.704
R1097 dvss.n415 dvss.n398 127.703
R1098 dvss.n547 dvss.n356 126.495
R1099 dvss.n511 dvss.n363 126.495
R1100 dvss.n609 dvss.t318 126.322
R1101 dvss.n596 dvss.t55 126.32
R1102 dvss.n457 dvss.n366 124.909
R1103 dvss.n162 dvss.t65 124.697
R1104 dvss.n297 dvss.t22 124.695
R1105 dvss.n1361 dvss.n1360 123.984
R1106 dvss.n1037 dvss.n1036 123.346
R1107 dvss.t410 dvss.t35 122.281
R1108 dvss.n766 dvss.t376 120.689
R1109 dvss.n766 dvss.t125 120.689
R1110 dvss.t81 dvss.t126 120.487
R1111 dvss.n950 dvss.n949 120.472
R1112 dvss.n413 dvss.n411 120.088
R1113 dvss.n1014 dvss.n930 119.806
R1114 dvss.n1030 dvss.n1028 119.575
R1115 dvss.n1054 dvss.n1053 118.722
R1116 dvss.n972 dvss.n971 117.001
R1117 dvss.n971 dvss.n789 117.001
R1118 dvss.n977 dvss.n963 117.001
R1119 dvss.n977 dvss.n976 117.001
R1120 dvss.n983 dvss.n931 117.001
R1121 dvss.n964 dvss.n931 117.001
R1122 dvss.n1013 dvss.n925 117.001
R1123 dvss.n1014 dvss.n1013 117.001
R1124 dvss.n1046 dvss.n1045 117.001
R1125 dvss.n1047 dvss.n1046 117.001
R1126 dvss.n1042 dvss.n1041 117.001
R1127 dvss.n1041 dvss.n1040 117.001
R1128 dvss.n1071 dvss.n852 117.001
R1129 dvss.n1082 dvss.n852 117.001
R1130 dvss.n1084 dvss.n1083 117.001
R1131 dvss.n1083 dvss.n1082 117.001
R1132 dvss.n846 dvss.n843 117.001
R1133 dvss.n846 dvss.n845 117.001
R1134 dvss.n1086 dvss.n1085 117.001
R1135 dvss.n1086 dvss.n845 117.001
R1136 dvss.n1030 dvss.n1029 117.001
R1137 dvss.n1029 dvss.n920 117.001
R1138 dvss.n1033 dvss.n1032 117.001
R1139 dvss.n1034 dvss.n1033 117.001
R1140 dvss.n932 dvss.n924 117.001
R1141 dvss.n932 dvss.n907 117.001
R1142 dvss.n1008 dvss.n1007 117.001
R1143 dvss.n1007 dvss.n1006 117.001
R1144 dvss.n955 dvss.n953 117.001
R1145 dvss.n955 dvss.n820 117.001
R1146 dvss.n951 dvss.n819 117.001
R1147 dvss.n1123 dvss.n819 117.001
R1148 dvss.n957 dvss.n956 117.001
R1149 dvss.n957 dvss.n820 117.001
R1150 dvss.n1125 dvss.n1124 117.001
R1151 dvss.n1124 dvss.n1123 117.001
R1152 dvss.n23 dvss.n22 117.001
R1153 dvss.n1418 dvss.n22 117.001
R1154 dvss.n1427 dvss.n1426 117.001
R1155 dvss.n1426 dvss.n1425 117.001
R1156 dvss.n1424 dvss.n1423 117.001
R1157 dvss.n1425 dvss.n1424 117.001
R1158 dvss.n1417 dvss.n21 117.001
R1159 dvss.n1418 dvss.n1417 117.001
R1160 dvss.n1301 dvss.n1300 117.001
R1161 dvss.t377 dvss.n1301 117.001
R1162 dvss.n1303 dvss.n1302 117.001
R1163 dvss.n1302 dvss.t377 117.001
R1164 dvss.n71 dvss.n69 117.001
R1165 dvss.n69 dvss.t237 117.001
R1166 dvss.n74 dvss.n70 117.001
R1167 dvss.n70 dvss.t237 117.001
R1168 dvss.n746 dvss.n741 117.001
R1169 dvss.n741 dvss.n738 117.001
R1170 dvss.n768 dvss.n767 117.001
R1171 dvss.n767 dvss.n766 117.001
R1172 dvss.n765 dvss.n764 117.001
R1173 dvss.n766 dvss.n765 117.001
R1174 dvss.n743 dvss.n740 117.001
R1175 dvss.n740 dvss.n738 117.001
R1176 dvss.n744 dvss.n739 117.001
R1177 dvss.n756 dvss.n739 117.001
R1178 dvss.n758 dvss.n757 117.001
R1179 dvss.n757 dvss.n756 117.001
R1180 dvss.t166 dvss.t83 114.403
R1181 dvss.t160 dvss.t420 113.793
R1182 dvss.n542 dvss.n362 113.695
R1183 dvss.n542 dvss.n541 113.695
R1184 dvss.n541 dvss.n540 113.695
R1185 dvss.n414 dvss.n413 113.695
R1186 dvss.n427 dvss.n414 113.695
R1187 dvss.n427 dvss.n426 113.695
R1188 dvss.n426 dvss.n415 113.695
R1189 dvss.t365 dvss.n738 112.507
R1190 dvss.n785 dvss.t248 112.233
R1191 dvss.n787 dvss.t63 112.233
R1192 dvss.t263 dvss.n638 111.538
R1193 dvss.n747 dvss.n746 110.438
R1194 dvss.t79 dvss.t75 109.632
R1195 dvss.n903 dvss.n887 108.906
R1196 dvss.n1377 dvss 108.642
R1197 dvss.n270 dvss.t134 108.198
R1198 dvss.t25 dvss.n245 108.198
R1199 dvss.n1147 dvss.n1146 107.272
R1200 dvss.n1386 dvss.t320 106.559
R1201 dvss.t322 dvss.n1386 106.559
R1202 dvss.n809 dvss.n808 105.412
R1203 dvss.n303 dvss.t21 104.486
R1204 dvss.n352 dvss.t14 104.486
R1205 dvss.n414 dvss.n410 103.906
R1206 dvss.n426 dvss.n425 103.906
R1207 dvss.n914 dvss.n913 103.906
R1208 dvss.n1109 dvss.n1108 103.906
R1209 dvss.n865 dvss.n848 103.772
R1210 dvss.n552 dvss.t90 103.306
R1211 dvss.n866 dvss.n865 101.944
R1212 dvss.n410 dvss.n400 101.647
R1213 dvss.n425 dvss.n401 101.647
R1214 dvss.t30 dvss.n456 101.198
R1215 dvss.n913 dvss.n825 100.141
R1216 dvss.n1109 dvss.n826 100.141
R1217 dvss.n239 dvss.n238 100.052
R1218 dvss.n230 dvss.n229 100.052
R1219 dvss.n216 dvss.n215 100.052
R1220 dvss.n209 dvss.n208 100.052
R1221 dvss.n198 dvss.n197 100.052
R1222 dvss.n185 dvss.n184 100.052
R1223 dvss.n172 dvss.n171 100.052
R1224 dvss.n582 dvss.n581 100.05
R1225 dvss.n576 dvss.n124 100.05
R1226 dvss.n560 dvss.n132 100.05
R1227 dvss.n346 dvss.n139 100.05
R1228 dvss.n332 dvss.n331 100.05
R1229 dvss.n326 dvss.n146 100.05
R1230 dvss.n310 dvss.n154 100.05
R1231 dvss.n521 dvss.n49 99.5749
R1232 dvss.n552 dvss.t226 99.0901
R1233 dvss.n500 dvss.t370 98.1874
R1234 dvss.n500 dvss.t109 98.1874
R1235 dvss.n731 dvss.t77 98.1874
R1236 dvss.n731 dvss.t205 98.1874
R1237 dvss.n756 dvss.n755 98.1874
R1238 dvss.t111 dvss.t340 98.1749
R1239 dvss.n540 dvss.n539 97.5005
R1240 dvss.n539 dvss.n538 97.5005
R1241 dvss.n543 dvss.n542 97.5005
R1242 dvss.n544 dvss.n543 97.5005
R1243 dvss.n513 dvss.n512 97.5005
R1244 dvss.n538 dvss.n513 97.5005
R1245 dvss.n546 dvss.n545 97.5005
R1246 dvss.n545 dvss.n544 97.5005
R1247 dvss.n918 dvss.n917 97.5005
R1248 dvss.n919 dvss.n918 97.5005
R1249 dvss.n913 dvss.n912 97.5005
R1250 dvss.n912 dvss.n829 97.5005
R1251 dvss.n1110 dvss.n1109 97.5005
R1252 dvss.n1111 dvss.n1110 97.5005
R1253 dvss.n1105 dvss.n834 97.5005
R1254 dvss.n1105 dvss.n1104 97.5005
R1255 dvss.n800 dvss.n795 97.5005
R1256 dvss.n800 dvss.n799 97.5005
R1257 dvss.n810 dvss.n798 97.5005
R1258 dvss.n1137 dvss.n798 97.5005
R1259 dvss.n1144 dvss.n1143 97.5005
R1260 dvss.n1145 dvss.n1144 97.5005
R1261 dvss.n76 dvss.n75 97.5005
R1262 dvss.n77 dvss.n76 97.5005
R1263 dvss.n73 dvss.n72 97.5005
R1264 dvss.n72 dvss.n27 97.5005
R1265 dvss.n421 dvss.n415 97.5005
R1266 dvss.n422 dvss.n421 97.5005
R1267 dvss.n428 dvss.n427 97.5005
R1268 dvss.n429 dvss.n428 97.5005
R1269 dvss.n413 dvss.n412 97.5005
R1270 dvss.n412 dvss.n367 97.5005
R1271 dvss.n411 dvss.n366 97.5005
R1272 dvss.n410 dvss.n409 97.5005
R1273 dvss.n409 dvss.n408 97.5005
R1274 dvss.n425 dvss.n424 97.5005
R1275 dvss.n424 dvss.n423 97.5005
R1276 dvss.n420 dvss.n418 97.5005
R1277 dvss.n420 dvss.n419 97.5005
R1278 dvss.n417 dvss.n416 97.5005
R1279 dvss.n422 dvss.n416 97.5005
R1280 dvss.n431 dvss.n430 97.5005
R1281 dvss.n430 dvss.n429 97.5005
R1282 dvss.n403 dvss.n402 97.5005
R1283 dvss.n403 dvss.n367 97.5005
R1284 dvss.n1072 dvss.n843 97.4474
R1285 dvss.n1092 dvss.n843 96.377
R1286 dvss.n930 dvss.n894 95.8456
R1287 dvss.n1300 dvss.n64 95.2476
R1288 dvss.n1300 dvss.n1299 95.2476
R1289 dvss.n926 dvss.n891 92.9825
R1290 dvss.n24 dvss.n21 92.4525
R1291 dvss.n639 dvss.t430 92.3082
R1292 dvss.n769 dvss.n82 91.8104
R1293 dvss.n651 dvss.n644 90.905
R1294 dvss.n1406 dvss.n1405 90.4228
R1295 dvss.n985 dvss.n962 89.1641
R1296 dvss.n1028 dvss.n903 88.375
R1297 dvss.n1130 dvss.n814 87.9969
R1298 dvss.n953 dvss.n952 87.9489
R1299 dvss.n652 dvss.n643 87.6306
R1300 dvss.n759 dvss.n758 87.3417
R1301 dvss.n1428 dvss.n1427 87.3417
R1302 dvss.n1427 dvss.n18 87.3417
R1303 dvss.n23 dvss.n18 87.3417
R1304 dvss.t419 dvss.t81 87.0188
R1305 dvss.t126 dvss.t60 87.0188
R1306 dvss.n503 dvss.n101 86.4507
R1307 dvss.n810 dvss.n809 85.4292
R1308 dvss.n570 dvss.t130 85.3191
R1309 dvss.n948 dvss.n946 84.8377
R1310 dvss.n915 dvss.n914 83.9534
R1311 dvss.n914 dvss.n833 83.9534
R1312 dvss.n1108 dvss.n833 83.9534
R1313 dvss.n1108 dvss.n1107 83.9534
R1314 dvss.n1155 dvss.n1149 83.7224
R1315 dvss.n989 dvss.n988 83.407
R1316 dvss.n986 dvss.n984 81.6649
R1317 dvss.n320 dvss.t138 81.267
R1318 dvss.n875 dvss.n872 81.2016
R1319 dvss.n1003 dvss.n935 80.6409
R1320 dvss.t32 dvss.t236 80.325
R1321 dvss.t236 dvss.t112 80.325
R1322 dvss.n362 dvss.n355 80.1887
R1323 dvss.t187 dvss.t410 80.1155
R1324 dvss.n533 dvss.n532 79.57
R1325 dvss.n524 dvss.n517 79.57
R1326 dvss.n502 dvss.n97 79.0593
R1327 dvss.n733 dvss.n97 79.0593
R1328 dvss.n734 dvss.n733 79.0593
R1329 dvss.n1392 dvss.n1381 79.0593
R1330 dvss.n1015 dvss.n1014 78.984
R1331 dvss.n373 dvss.t386 76.8564
R1332 dvss.n1295 dvss.n1294 75.8227
R1333 dvss.n973 dvss.n972 75.4543
R1334 dvss.n419 dvss.t46 73.7906
R1335 dvss.n554 dvss.n553 73.5273
R1336 dvss.n745 dvss.n736 73.0738
R1337 dvss.n747 dvss.n745 72.206
R1338 dvss.n1165 dvss.t338 71.9283
R1339 dvss.n1162 dvss.t39 71.9283
R1340 dvss.n529 dvss.n518 71.5299
R1341 dvss.n759 dvss.n735 71.5299
R1342 dvss.n742 dvss.n735 71.5299
R1343 dvss.n734 dvss.n96 71.5299
R1344 dvss.n96 dvss.n87 71.5299
R1345 dvss.n100 dvss.n97 71.5299
R1346 dvss.n724 dvss.n100 71.5299
R1347 dvss.n725 dvss.n82 71.5299
R1348 dvss.n91 dvss.n88 71.5299
R1349 dvss.n91 dvss.n83 71.5299
R1350 dvss.n17 dvss.n6 71.5299
R1351 dvss.n1428 dvss.n17 71.5299
R1352 dvss.n14 dvss.n5 71.5299
R1353 dvss.n15 dvss.n14 71.5299
R1354 dvss.n1394 dvss.n1383 71.5299
R1355 dvss.n1399 dvss.n1394 71.5299
R1356 dvss.n1404 dvss.n1382 71.5299
R1357 dvss.n1392 dvss.n1382 71.5299
R1358 dvss.n1422 dvss.n1421 71.5299
R1359 dvss.n1421 dvss.n18 71.5299
R1360 dvss.n1065 dvss.n867 71.2831
R1361 dvss.n530 dvss.n529 70.777
R1362 dvss.n1006 dvss.n937 70.1793
R1363 dvss.n1019 dvss.n1018 70.0532
R1364 dvss.n1017 dvss.n891 69.1602
R1365 dvss.n438 dvss.n437 68.8522
R1366 dvss.n438 dvss.n436 68.7355
R1367 dvss.n439 dvss.n435 68.7333
R1368 dvss.n973 dvss.n963 66.6531
R1369 dvss.n418 dvss.n417 66.3047
R1370 dvss.n1044 dvss.n901 65.9625
R1371 dvss.n1003 dvss.n1002 65.4191
R1372 dvss.n456 dvss.n367 65.3575
R1373 dvss.n1052 dvss.n890 65.1217
R1374 dvss.n508 dvss.n363 65.0005
R1375 dvss.n509 dvss.n508 65.0005
R1376 dvss.n365 dvss.n364 65.0005
R1377 dvss.n537 dvss.n365 65.0005
R1378 dvss.n550 dvss.n549 65.0005
R1379 dvss.n551 dvss.n550 65.0005
R1380 dvss.n372 dvss.n356 65.0005
R1381 dvss.n373 dvss.n372 65.0005
R1382 dvss.n1094 dvss.n838 65.0005
R1383 dvss.n883 dvss.n838 65.0005
R1384 dvss.n1075 dvss.n849 65.0005
R1385 dvss.n851 dvss.n849 65.0005
R1386 dvss.n1077 dvss.n850 65.0005
R1387 dvss.n1081 dvss.n850 65.0005
R1388 dvss.n841 dvss.n839 65.0005
R1389 dvss.n839 dvss.n837 65.0005
R1390 dvss.n1307 dvss.n1306 65.0005
R1391 dvss.n1308 dvss.n1307 65.0005
R1392 dvss.n61 dvss.n54 65.0005
R1393 dvss.n61 dvss.n59 65.0005
R1394 dvss.n66 dvss.n65 65.0005
R1395 dvss.n65 dvss.n60 65.0005
R1396 dvss.n68 dvss.n67 65.0005
R1397 dvss.n78 dvss.n68 65.0005
R1398 dvss.t374 dvss.n192 64.9185
R1399 dvss.n604 dvss.t317 64.9185
R1400 dvss.n916 dvss.n825 64.8732
R1401 dvss.n1114 dvss.n826 64.8732
R1402 dvss.n835 dvss.n826 64.8732
R1403 dvss.n1115 dvss.n825 64.2914
R1404 dvss.n1312 dvss.t412 63.375
R1405 dvss.n616 dvss.t259 62.8576
R1406 dvss.n1134 dvss.n804 62.758
R1407 dvss.n808 dvss.n794 62.4946
R1408 dvss.n1347 dvss.t84 62.2404
R1409 dvss.n1058 dvss.n887 61.5624
R1410 dvss.n587 dvss.t70 60.9423
R1411 dvss.n402 dvss.n399 60.3224
R1412 dvss.t61 dvss.n1313 60.2439
R1413 dvss.n967 dvss.n966 60.2175
R1414 dvss.n518 dvss.n516 59.4829
R1415 dvss.n525 dvss.n518 59.4829
R1416 dvss.n760 dvss.n734 59.4829
R1417 dvss.n760 dvss.n759 59.4829
R1418 dvss.n1400 dvss.n1392 59.4829
R1419 dvss.n1400 dvss.n1399 59.4829
R1420 dvss.n1399 dvss.n1398 59.4829
R1421 dvss.n1398 dvss.n15 59.4829
R1422 dvss.n1429 dvss.n15 59.4829
R1423 dvss.n1429 dvss.n1428 59.4829
R1424 dvss.n1094 dvss.n1093 59.2721
R1425 dvss.n1334 dvss.t33 59.2552
R1426 dvss.n337 dvss.t92 58.048
R1427 dvss.t83 dvss.n1312 55.9188
R1428 dvss.n42 dvss.t82 55.7148
R1429 dvss.n42 dvss.t127 55.7148
R1430 dvss.n905 dvss.n897 51.4729
R1431 dvss.n1305 dvss.n1304 50.6672
R1432 dvss.t185 dvss.t121 50.5994
R1433 dvss.n689 dvss.t261 49.8075
R1434 dvss.n441 dvss.t159 49.3953
R1435 dvss.n1048 dvss.n1047 48.8105
R1436 dvss.n974 dvss.n973 48.7505
R1437 dvss.n975 dvss.n974 48.7505
R1438 dvss.n979 dvss.n978 48.7505
R1439 dvss.n1093 dvss.n1092 48.0896
R1440 dvss.n45 dvss.t421 47.6797
R1441 dvss.n1360 dvss.t6 47.2956
R1442 dvss.n981 dvss.n980 46.2264
R1443 dvss.n408 dvss.t42 44.2746
R1444 dvss.t35 dvss.n422 44.2746
R1445 dvss.n1292 dvss.t209 43.6661
R1446 dvss.n1143 dvss.n1142 43.5408
R1447 dvss.n729 dvss.t376 42.9573
R1448 dvss.n775 dvss.t378 42.478
R1449 dvss.n1064 dvss.n1063 41.7862
R1450 dvss.n1063 dvss.n1062 41.7862
R1451 dvss.n880 dvss.n879 41.7862
R1452 dvss.n881 dvss.n880 41.7862
R1453 dvss.n53 dvss.n51 41.7862
R1454 dvss.n58 dvss.n51 41.7862
R1455 dvss.n1305 dvss.n52 41.7862
R1456 dvss.n58 dvss.n52 41.7862
R1457 dvss.n982 dvss.n981 41.5158
R1458 dvss.n873 dvss.n868 41.5006
R1459 dvss.n689 dvss.t431 41.3519
R1460 dvss.n984 dvss.n982 41.2882
R1461 dvss.n988 dvss.n961 40.465
R1462 dvss.n397 dvss.n396 40.2093
R1463 dvss.n712 dvss.n105 40.2093
R1464 dvss.n616 dvss.t74 40.0005
R1465 dvss.n395 dvss.t391 39.6005
R1466 dvss.n395 dvss.t215 39.6005
R1467 dvss.n394 dvss.t200 39.6005
R1468 dvss.n394 dvss.t439 39.6005
R1469 dvss.n393 dvss.t221 39.6005
R1470 dvss.n393 dvss.t393 39.6005
R1471 dvss.n392 dvss.t227 39.6005
R1472 dvss.n392 dvss.t91 39.6005
R1473 dvss.n391 dvss.t41 39.6005
R1474 dvss.n391 dvss.t241 39.6005
R1475 dvss.n390 dvss.t169 39.6005
R1476 dvss.n390 dvss.t47 39.6005
R1477 dvss.n378 dvss.t36 39.6005
R1478 dvss.n378 dvss.t211 39.6005
R1479 dvss.n379 dvss.t105 39.6005
R1480 dvss.n379 dvss.t188 39.6005
R1481 dvss.n380 dvss.t192 39.6005
R1482 dvss.n380 dvss.t382 39.6005
R1483 dvss.n381 dvss.t306 39.6005
R1484 dvss.n381 dvss.t186 39.6005
R1485 dvss.n382 dvss.t101 39.6005
R1486 dvss.n382 dvss.t190 39.6005
R1487 dvss.n383 dvss.t103 39.6005
R1488 dvss.n383 dvss.t43 39.6005
R1489 dvss.n443 dvss.t213 39.6005
R1490 dvss.n443 dvss.t387 39.6005
R1491 dvss.n472 dvss.t97 39.6005
R1492 dvss.n472 dvss.t165 39.6005
R1493 dvss.n471 dvss.t231 39.6005
R1494 dvss.n471 dvss.t406 39.6005
R1495 dvss.n470 dvss.t99 39.6005
R1496 dvss.n470 dvss.t233 39.6005
R1497 dvss.n469 dvss.t302 39.6005
R1498 dvss.n469 dvss.t308 39.6005
R1499 dvss.n468 dvss.t385 39.6005
R1500 dvss.n468 dvss.t434 39.6005
R1501 dvss.n467 dvss.t404 39.6005
R1502 dvss.n467 dvss.t300 39.6005
R1503 dvss.n479 dvss.t120 39.6005
R1504 dvss.n479 dvss.t163 39.6005
R1505 dvss.n480 dvss.t304 39.6005
R1506 dvss.n480 dvss.t268 39.6005
R1507 dvss.n481 dvss.t57 39.6005
R1508 dvss.n481 dvss.t278 39.6005
R1509 dvss.n482 dvss.t270 39.6005
R1510 dvss.n482 dvss.t274 39.6005
R1511 dvss.n483 dvss.t59 39.6005
R1512 dvss.n483 dvss.t272 39.6005
R1513 dvss.n484 dvss.t276 39.6005
R1514 dvss.n484 dvss.t337 39.6005
R1515 dvss.n102 dvss.t335 39.6005
R1516 dvss.n102 dvss.t235 39.6005
R1517 dvss.n0 dvss.t321 39.6005
R1518 dvss.n0 dvss.t323 39.6005
R1519 dvss.n1079 dvss.n1078 39.0005
R1520 dvss.n1080 dvss.n1079 39.0005
R1521 dvss.n877 dvss.n876 39.0005
R1522 dvss.n876 dvss.n871 39.0005
R1523 dvss.n1132 dvss.n1131 39.0005
R1524 dvss.n1133 dvss.n1132 39.0005
R1525 dvss.n948 dvss.n947 39.0005
R1526 dvss.n947 dvss.n803 39.0005
R1527 dvss.n954 dvss.n942 39.0005
R1528 dvss.n944 dvss.n942 39.0005
R1529 dvss.n996 dvss.n940 39.0005
R1530 dvss.n997 dvss.n996 39.0005
R1531 dvss.n1004 dvss.n1003 39.0005
R1532 dvss.n1005 dvss.n1004 39.0005
R1533 dvss.t203 dvss.t125 38.8661
R1534 dvss.n768 dvss.n83 38.5667
R1535 dvss.n746 dvss.n83 38.5667
R1536 dvss.n987 dvss.n962 38.4005
R1537 dvss.n589 dvss.t54 36.5656
R1538 dvss.n707 dvss.n614 36.1417
R1539 dvss.n702 dvss.n701 36.1417
R1540 dvss.n697 dvss.n696 36.1417
R1541 dvss.n696 dvss.n695 36.1417
R1542 dvss.n695 dvss.n619 36.1417
R1543 dvss.n691 dvss.n619 36.1417
R1544 dvss.n687 dvss.n621 36.1417
R1545 dvss.n683 dvss.n621 36.1417
R1546 dvss.n683 dvss.n682 36.1417
R1547 dvss.n682 dvss.n681 36.1417
R1548 dvss.n675 dvss.n626 36.1417
R1549 dvss.n664 dvss.n663 36.1417
R1550 dvss.n1321 dvss.n1320 36.1417
R1551 dvss.n1322 dvss.n1321 36.1417
R1552 dvss.n1327 dvss.n1326 36.1417
R1553 dvss.n1328 dvss.n1327 36.1417
R1554 dvss.n1328 dvss.n40 36.1417
R1555 dvss.n1332 dvss.n40 36.1417
R1556 dvss.n1333 dvss.n1332 36.1417
R1557 dvss.n1339 dvss.n38 36.1417
R1558 dvss.n1340 dvss.n1339 36.1417
R1559 dvss.n1341 dvss.n1340 36.1417
R1560 dvss.n1341 dvss.n36 36.1417
R1561 dvss.n1352 dvss.n34 36.1417
R1562 dvss.n1353 dvss.n1352 36.1417
R1563 dvss.n1355 dvss.n32 36.1417
R1564 dvss.n1359 dvss.n32 36.1417
R1565 dvss.n1363 dvss.n1362 36.1417
R1566 dvss.n290 dvss.n289 36.1417
R1567 dvss.n289 dvss.n288 36.1417
R1568 dvss.n288 dvss.n165 36.1417
R1569 dvss.n282 dvss.n165 36.1417
R1570 dvss.n282 dvss.n281 36.1417
R1571 dvss.n281 dvss.n280 36.1417
R1572 dvss.n280 dvss.n176 36.1417
R1573 dvss.n274 dvss.n176 36.1417
R1574 dvss.n274 dvss.n273 36.1417
R1575 dvss.n273 dvss.n272 36.1417
R1576 dvss.n272 dvss.n189 36.1417
R1577 dvss.n266 dvss.n189 36.1417
R1578 dvss.n266 dvss.n265 36.1417
R1579 dvss.n265 dvss.n264 36.1417
R1580 dvss.n264 dvss.n203 36.1417
R1581 dvss.n258 dvss.n203 36.1417
R1582 dvss.n258 dvss.n257 36.1417
R1583 dvss.n257 dvss.n256 36.1417
R1584 dvss.n256 dvss.n219 36.1417
R1585 dvss.n250 dvss.n219 36.1417
R1586 dvss.n250 dvss.n249 36.1417
R1587 dvss.n249 dvss.n248 36.1417
R1588 dvss.n248 dvss.n233 36.1417
R1589 dvss.n242 dvss.n233 36.1417
R1590 dvss.n242 dvss.n111 36.1417
R1591 dvss.n606 dvss.n111 36.1417
R1592 dvss.n606 dvss.n112 36.1417
R1593 dvss.n300 dvss.n295 36.1417
R1594 dvss.n300 dvss.n156 36.1417
R1595 dvss.n307 dvss.n156 36.1417
R1596 dvss.n307 dvss.n152 36.1417
R1597 dvss.n314 dvss.n152 36.1417
R1598 dvss.n314 dvss.n148 36.1417
R1599 dvss.n323 dvss.n148 36.1417
R1600 dvss.n323 dvss.n322 36.1417
R1601 dvss.n322 dvss.n144 36.1417
R1602 dvss.n335 dvss.n144 36.1417
R1603 dvss.n335 dvss.n141 36.1417
R1604 dvss.n342 dvss.n141 36.1417
R1605 dvss.n342 dvss.n137 36.1417
R1606 dvss.n349 dvss.n137 36.1417
R1607 dvss.n349 dvss.n134 36.1417
R1608 dvss.n557 dvss.n134 36.1417
R1609 dvss.n557 dvss.n130 36.1417
R1610 dvss.n564 dvss.n130 36.1417
R1611 dvss.n564 dvss.n126 36.1417
R1612 dvss.n573 dvss.n126 36.1417
R1613 dvss.n573 dvss.n572 36.1417
R1614 dvss.n572 dvss.n122 36.1417
R1615 dvss.n585 dvss.n122 36.1417
R1616 dvss.n585 dvss.n119 36.1417
R1617 dvss.n592 dvss.n119 36.1417
R1618 dvss.n592 dvss.n117 36.1417
R1619 dvss.n599 dvss.n117 36.1417
R1620 dvss.n1049 dvss.n894 35.4987
R1621 dvss.n1290 dvss.n777 35.4084
R1622 dvss.n1291 dvss.n776 35.4054
R1623 dvss.n773 dvss.n80 35.4029
R1624 dvss.n1289 dvss.n778 35.3969
R1625 dvss.n774 dvss.n79 35.3787
R1626 dvss.n1335 dvss.n38 35.0123
R1627 dvss.n339 dvss.t293 34.829
R1628 dvss.n1150 dvss.t429 34.8005
R1629 dvss.n1150 dvss.t427 34.8005
R1630 dvss.n1151 dvss.t399 34.8005
R1631 dvss.n1151 dvss.t402 34.8005
R1632 dvss.n1011 dvss.n1010 34.4123
R1633 dvss.n1011 dvss.n929 34.4123
R1634 dvss.n1026 dvss.n1025 34.4123
R1635 dvss.n1025 dvss.n894 34.4123
R1636 dvss.n922 dvss.n902 34.4123
R1637 dvss.n922 dvss.n905 34.4123
R1638 dvss.n1028 dvss.n904 34.4123
R1639 dvss.n1039 dvss.n904 34.4123
R1640 dvss.n985 dvss.n936 34.4123
R1641 dvss.n965 dvss.n936 34.4123
R1642 dvss.n628 dvss.t144 34.0546
R1643 dvss.n628 dvss.t156 34.0546
R1644 dvss.n630 dvss.t150 34.0546
R1645 dvss.n630 dvss.t148 34.0546
R1646 dvss.n633 dvss.t154 34.0546
R1647 dvss.n961 dvss.n960 33.6801
R1648 dvss.n668 dvss.n631 33.1299
R1649 dvss.n1087 dvss.n844 32.5005
R1650 dvss.n1088 dvss.n1087 32.5005
R1651 dvss.n1073 dvss.n847 32.5005
R1652 dvss.n1036 dvss.n847 32.5005
R1653 dvss.n1121 dvss.n1120 32.5005
R1654 dvss.n1122 dvss.n1121 32.5005
R1655 dvss.n817 dvss.n813 32.5005
R1656 dvss.n817 dvss.n805 32.5005
R1657 dvss.n960 dvss.n959 32.5005
R1658 dvss.n959 dvss.n958 32.5005
R1659 dvss.n623 dvss.t254 32.4329
R1660 dvss.n623 dvss.t8 32.4329
R1661 dvss.n952 dvss.n822 32.3833
R1662 dvss.t158 dvss.t214 32.0238
R1663 dvss.n1363 dvss.n30 32.0005
R1664 dvss.n402 dvss.n400 31.6857
R1665 dvss.n431 dvss.n401 31.6857
R1666 dvss.n417 dvss.n401 31.6857
R1667 dvss.n703 dvss.n614 31.2476
R1668 dvss.n1054 dvss.n1052 30.8082
R1669 dvss.n992 dvss.n935 30.6755
R1670 dvss.n1119 dvss.n816 30.1319
R1671 dvss.n677 dvss.n676 30.1181
R1672 dvss.n670 dvss.n669 30.1181
R1673 dvss.n688 dvss.n687 30.0632
R1674 dvss.n637 dvss.t289 30.0005
R1675 dvss.n868 dvss.n867 29.7851
R1676 dvss.n432 dvss.n400 29.5874
R1677 dvss.n1316 dvss.n46 29.3652
R1678 dvss.n954 dvss.n941 29.3251
R1679 dvss.n1168 dvss.n780 29.3166
R1680 dvss.n1345 dvss.n36 28.9887
R1681 dvss.n1348 dvss.n1346 28.9887
R1682 dvss.n677 dvss.n624 28.6123
R1683 dvss.n662 dvss.n635 28.6123
R1684 dvss.n1009 dvss.n1008 27.7719
R1685 dvss.n1009 dvss.n924 27.7719
R1686 dvss.n1027 dvss.n924 27.7719
R1687 dvss.n1032 dvss.n1027 27.7719
R1688 dvss.n1032 dvss.n1031 27.7719
R1689 dvss.n1031 dvss.n1030 27.7719
R1690 dvss.n1091 dvss.n844 26.9228
R1691 dvss.n708 dvss.n707 26.7299
R1692 dvss.n671 dvss.n626 26.7299
R1693 dvss.n1374 dvss.n1369 25.977
R1694 dvss.n970 dvss.n969 25.7896
R1695 dvss.n1346 dvss.n1345 25.6005
R1696 dvss.n980 dvss.n979 25.2546
R1697 dvss.n656 dvss.n641 24.8476
R1698 dvss.n1316 dvss.n1315 24.8476
R1699 dvss.n1376 dvss.n1375 24.8476
R1700 dvss.n966 dvss.n788 24.6159
R1701 dvss.n1120 dvss.n1119 24.4927
R1702 dvss.n701 dvss.n617 24.4711
R1703 dvss.n658 dvss.n657 24.4711
R1704 dvss.n1322 dvss.n43 24.4711
R1705 dvss.n1348 dvss.n34 24.4711
R1706 dvss.n1298 dvss.n1297 24.3755
R1707 dvss.n1297 dvss.t228 24.3755
R1708 dvss.n1296 dvss.n1295 24.3755
R1709 dvss.t228 dvss.n1296 24.3755
R1710 dvss.n991 dvss.n990 24.2648
R1711 dvss.n1320 dvss.n46 24.0946
R1712 dvss.n979 dvss.n970 23.914
R1713 dvss.n676 dvss.n675 23.3417
R1714 dvss.n697 dvss.n617 22.9652
R1715 dvss.n657 dvss.n656 22.9652
R1716 dvss.n1347 dvss.t167 22.7037
R1717 dvss.n633 dvss.t146 22.7032
R1718 dvss.n634 dvss.t152 22.7032
R1719 dvss.n634 dvss.t287 22.7032
R1720 dvss.n637 dvss.t285 22.7032
R1721 dvss.n1304 dvss.n1303 22.4894
R1722 dvss.n1303 dvss.n55 22.4894
R1723 dvss.n808 dvss.n795 22.3548
R1724 dvss.n1282 dvss.n1253 22.3023
R1725 dvss.n703 dvss.n702 22.2123
R1726 dvss.n972 dvss.n970 22.2123
R1727 dvss.n969 dvss.n889 22.0715
R1728 dvss.n877 dvss.n875 22.0326
R1729 dvss.n1360 dvss.t281 21.9347
R1730 dvss.n810 dvss.n796 21.7696
R1731 dvss.n178 dvss.t309 21.6398
R1732 dvss.n254 dvss.t313 21.6398
R1733 dvss.n1141 dvss.n795 21.5764
R1734 dvss.n779 dvss.t246 21.5736
R1735 dvss.n45 dvss.t161 21.551
R1736 dvss.n1065 dvss.n1064 21.4672
R1737 dvss.n238 dvss.t26 21.2805
R1738 dvss.n238 dvss.t24 21.2805
R1739 dvss.n229 dvss.t67 21.2805
R1740 dvss.n229 dvss.t17 21.2805
R1741 dvss.n215 dvss.t69 21.2805
R1742 dvss.n215 dvss.t314 21.2805
R1743 dvss.n208 dvss.t375 21.2805
R1744 dvss.n208 dvss.t137 21.2805
R1745 dvss.n197 dvss.t135 21.2805
R1746 dvss.n197 dvss.t87 21.2805
R1747 dvss.n184 dvss.t296 21.2805
R1748 dvss.n184 dvss.t95 21.2805
R1749 dvss.n171 dvss.t223 21.2805
R1750 dvss.n171 dvss.t310 21.2805
R1751 dvss.n581 dvss.t71 21.2805
R1752 dvss.n581 dvss.t129 21.2805
R1753 dvss.n124 dvss.t217 21.2805
R1754 dvss.n124 dvss.t131 21.2805
R1755 dvss.n132 dvss.t219 21.2805
R1756 dvss.n132 dvss.t1 21.2805
R1757 dvss.n139 dvss.t294 21.2805
R1758 dvss.n139 dvss.t15 21.2805
R1759 dvss.n331 dvss.t93 21.2805
R1760 dvss.n331 dvss.t312 21.2805
R1761 dvss.n146 dvss.t266 21.2805
R1762 dvss.n146 dvss.t139 21.2805
R1763 dvss.n154 dvss.t133 21.2805
R1764 dvss.n154 dvss.t373 21.2805
R1765 dvss.n1281 dvss.n1254 21.1647
R1766 dvss.n691 dvss.n690 21.1456
R1767 dvss.t189 dvss.t107 21.0834
R1768 dvss.n1267 dvss.n1261 20.8934
R1769 dvss.n1261 dvss.n1260 20.8934
R1770 dvss.n671 dvss.n670 20.7064
R1771 dvss.n1423 dvss.n6 20.4805
R1772 dvss.n1423 dvss.n1422 20.4805
R1773 dvss.n1422 dvss.n21 20.4805
R1774 dvss.t350 dvss.n750 20.4751
R1775 dvss.t205 dvss.n730 20.4561
R1776 dvss.n1376 dvss.n30 19.9534
R1777 dvss.n547 dvss.n546 19.2323
R1778 dvss.n512 dvss.n511 19.2323
R1779 dvss.n681 dvss.n624 18.824
R1780 dvss.n658 dvss.n635 18.824
R1781 dvss.n377 dvss.n376 18.6433
R1782 dvss.n494 dvss.n493 18.6433
R1783 dvss.n1405 dvss.n1404 18.5384
R1784 dvss.n769 dvss.n768 18.2862
R1785 dvss.n956 dvss.n941 18.1745
R1786 dvss.n669 dvss.n668 17.3181
R1787 dvss.n1091 dvss.n1090 17.2064
R1788 dvss.n1090 dvss.n1089 17.2064
R1789 dvss.n1102 dvss.n1101 17.2064
R1790 dvss.n1103 dvss.n1102 17.2064
R1791 dvss.n1375 dvss.n1374 16.9417
R1792 dvss.n437 dvss.t31 16.5305
R1793 dvss.n437 dvss.t76 16.5305
R1794 dvss.n436 dvss.t108 16.5305
R1795 dvss.n436 dvss.t122 16.5305
R1796 dvss.n435 dvss.t411 16.5305
R1797 dvss.n435 dvss.t244 16.5305
R1798 dvss.n982 dvss.n928 16.2505
R1799 dvss.n927 dvss.n926 16.2505
R1800 dvss.n1064 dvss.n868 16.1338
R1801 dvss.n1125 dvss.n816 15.7807
R1802 dvss.n1000 dvss.n941 15.7807
R1803 dvss.n1126 dvss.n814 15.4875
R1804 dvss.n1076 dvss.n1075 15.4479
R1805 dvss.n709 dvss.n708 15.4358
R1806 dvss.n980 dvss.n963 15.3345
R1807 dvss.n945 dvss.n814 15.0967
R1808 dvss.n462 dvss.n460 15.0005
R1809 dvss.t119 dvss.n460 15.0005
R1810 dvss.n461 dvss.n459 15.0005
R1811 dvss.t119 dvss.n459 15.0005
R1812 dvss.n371 dvss.n369 15.0005
R1813 dvss.t168 dvss.n369 15.0005
R1814 dvss.n370 dvss.n368 15.0005
R1815 dvss.t168 dvss.n368 15.0005
R1816 dvss.n1146 dvss.n788 14.7987
R1817 dvss.n1271 dvss.n1254 14.7701
R1818 dvss.n429 dvss.t305 14.7585
R1819 dvss.n423 dvss.t381 14.7585
R1820 dvss.n1326 dvss.n43 14.6829
R1821 dvss.n901 dvss.n893 14.6255
R1822 dvss.n1048 dvss.n893 14.6255
R1823 dvss.n1018 dvss.n892 14.6255
R1824 dvss.n930 dvss.n892 14.6255
R1825 dvss.n726 dvss.n724 14.5302
R1826 dvss.n743 dvss.n742 14.448
R1827 dvss.n745 dvss.n744 14.3554
R1828 dvss.n755 dvss.t201 14.3142
R1829 dvss.n664 dvss.n631 14.3064
R1830 dvss.n511 dvss.n357 14.1378
R1831 dvss.n1404 dvss.n1403 13.9481
R1832 dvss.n1403 dvss.n1383 13.9481
R1833 dvss.n1395 dvss.n1383 13.9481
R1834 dvss.n1395 dvss.n5 13.9481
R1835 dvss.n1432 dvss.n6 13.9481
R1836 dvss.n1141 dvss.n1140 13.6799
R1837 dvss.n1060 dvss.n1059 13.6052
R1838 dvss.n1061 dvss.n1060 13.6052
R1839 dvss.n969 dvss.n968 13.6052
R1840 dvss.n1017 dvss.n1016 13.6052
R1841 dvss.n1016 dvss.n1015 13.6052
R1842 dvss.n896 dvss.n890 13.6052
R1843 dvss.n897 dvss.n896 13.6052
R1844 dvss.n783 dvss.n781 13.6052
R1845 dvss.n787 dvss.n783 13.6052
R1846 dvss.n782 dvss.n780 13.6052
R1847 dvss.n782 dvss.n26 13.6052
R1848 dvss.n1159 dvss.n1148 13.6052
R1849 dvss.n1148 dvss.n1147 13.6052
R1850 dvss.n1156 dvss.n786 13.6052
R1851 dvss.n786 dvss.n785 13.6052
R1852 dvss.n548 dvss.n547 13.5647
R1853 dvss.n1078 dvss.n1077 13.5534
R1854 dvss.n723 dvss.n101 13.2848
R1855 dvss.n551 dvss.t438 12.8098
R1856 dvss.n1335 dvss.n1333 12.424
R1857 dvss.n1078 dvss.n856 12.1845
R1858 dvss.n872 dvss.n856 12.0414
R1859 dvss.n946 dvss.n945 11.9211
R1860 dvss.t372 dvss.n150 11.61
R1861 dvss.t0 dvss.n128 11.61
R1862 dvss.n875 dvss.n874 11.4592
R1863 dvss.n1369 dvss.n1368 11.4477
R1864 dvss.n1074 dvss.n1073 11.405
R1865 dvss.n663 dvss.n662 11.2946
R1866 dvss.n1052 dvss.n1051 11.2477
R1867 dvss.n1271 dvss.n1270 11.2225
R1868 dvss.n1051 dvss.n891 10.912
R1869 dvss.n1001 dvss.n1000 10.6509
R1870 dvss.n1002 dvss.n1001 10.6509
R1871 dvss.n1362 dvss.n1361 10.5417
R1872 dvss.n956 dvss.n816 10.4066
R1873 dvss.n946 dvss.n796 10.26
R1874 dvss.n753 dvss.t407 10.2283
R1875 dvss.n1092 dvss.n1091 10.1559
R1876 dvss.n763 dvss.n88 9.75892
R1877 dvss.n725 dvss.n87 9.63218
R1878 dvss.n887 dvss.n885 9.59066
R1879 dvss.n906 dvss.n885 9.59066
R1880 dvss.n1053 dvss.n884 9.59066
R1881 dvss.n906 dvss.n884 9.59066
R1882 dvss.n1130 dvss.n1129 9.35854
R1883 dvss.n1269 dvss.n1253 9.35596
R1884 dvss.n296 dvss.n295 9.34345
R1885 dvss.n290 dvss.n160 9.34253
R1886 dvss.n1315 dvss 9.3308
R1887 dvss.n1370 dvss.n1369 9.3005
R1888 dvss.n1317 dvss.n1316 9.3005
R1889 dvss.n1318 dvss.n46 9.3005
R1890 dvss.n1320 dvss.n1319 9.3005
R1891 dvss.n1321 dvss.n44 9.3005
R1892 dvss.n1323 dvss.n1322 9.3005
R1893 dvss.n1324 dvss.n43 9.3005
R1894 dvss.n1326 dvss.n1325 9.3005
R1895 dvss.n1327 dvss.n41 9.3005
R1896 dvss.n1329 dvss.n1328 9.3005
R1897 dvss.n1330 dvss.n40 9.3005
R1898 dvss.n1332 dvss.n1331 9.3005
R1899 dvss.n1333 dvss.n39 9.3005
R1900 dvss.n1336 dvss.n1335 9.3005
R1901 dvss.n1337 dvss.n38 9.3005
R1902 dvss.n1339 dvss.n1338 9.3005
R1903 dvss.n1340 dvss.n37 9.3005
R1904 dvss.n1342 dvss.n1341 9.3005
R1905 dvss.n1343 dvss.n36 9.3005
R1906 dvss.n1345 dvss.n1344 9.3005
R1907 dvss.n1346 dvss.n35 9.3005
R1908 dvss.n1349 dvss.n1348 9.3005
R1909 dvss.n1350 dvss.n34 9.3005
R1910 dvss.n1352 dvss.n1351 9.3005
R1911 dvss.n1353 dvss.n33 9.3005
R1912 dvss.n1356 dvss.n1355 9.3005
R1913 dvss.n1357 dvss.n32 9.3005
R1914 dvss.n1359 dvss.n1358 9.3005
R1915 dvss.n1362 dvss.n31 9.3005
R1916 dvss.n1364 dvss.n1363 9.3005
R1917 dvss.n1376 dvss.n1366 9.3005
R1918 dvss.n1375 dvss.n1367 9.3005
R1919 dvss.n1374 dvss.n1373 9.3005
R1920 dvss.n1372 dvss.n1369 9.3005
R1921 dvss.n163 dvss.n162 9.3005
R1922 dvss.n162 dvss.n160 9.3005
R1923 dvss.n172 dvss.n170 9.3005
R1924 dvss.n186 dvss.n185 9.3005
R1925 dvss.n185 dvss.n183 9.3005
R1926 dvss.n185 dvss.n181 9.3005
R1927 dvss.n199 dvss.n198 9.3005
R1928 dvss.n198 dvss.n196 9.3005
R1929 dvss.n198 dvss.n195 9.3005
R1930 dvss.n210 dvss.n209 9.3005
R1931 dvss.n209 dvss.n207 9.3005
R1932 dvss.n209 dvss.n206 9.3005
R1933 dvss.n216 dvss.n214 9.3005
R1934 dvss.n231 dvss.n230 9.3005
R1935 dvss.n230 dvss.n228 9.3005
R1936 dvss.n230 dvss.n227 9.3005
R1937 dvss.n240 dvss.n239 9.3005
R1938 dvss.n239 dvss.n235 9.3005
R1939 dvss.n239 dvss.n237 9.3005
R1940 dvss.n610 dvss.n609 9.3005
R1941 dvss.n609 dvss.n608 9.3005
R1942 dvss.n289 dvss.n161 9.3005
R1943 dvss.n288 dvss.n164 9.3005
R1944 dvss.n169 dvss.n165 9.3005
R1945 dvss.n282 dvss.n168 9.3005
R1946 dvss.n281 dvss.n174 9.3005
R1947 dvss.n280 dvss.n175 9.3005
R1948 dvss.n182 dvss.n176 9.3005
R1949 dvss.n274 dvss.n180 9.3005
R1950 dvss.n273 dvss.n187 9.3005
R1951 dvss.n272 dvss.n188 9.3005
R1952 dvss.n194 dvss.n189 9.3005
R1953 dvss.n266 dvss.n200 9.3005
R1954 dvss.n265 dvss.n201 9.3005
R1955 dvss.n264 dvss.n202 9.3005
R1956 dvss.n211 dvss.n203 9.3005
R1957 dvss.n258 dvss.n212 9.3005
R1958 dvss.n257 dvss.n213 9.3005
R1959 dvss.n256 dvss.n218 9.3005
R1960 dvss.n226 dvss.n219 9.3005
R1961 dvss.n250 dvss.n224 9.3005
R1962 dvss.n249 dvss.n225 9.3005
R1963 dvss.n248 dvss.n232 9.3005
R1964 dvss.n236 dvss.n233 9.3005
R1965 dvss.n242 dvss.n241 9.3005
R1966 dvss.n111 dvss.n110 9.3005
R1967 dvss.n607 dvss.n606 9.3005
R1968 dvss.n112 dvss.n109 9.3005
R1969 dvss.n298 dvss.n297 9.3005
R1970 dvss.n297 dvss.n296 9.3005
R1971 dvss.n310 dvss.n309 9.3005
R1972 dvss.n327 dvss.n326 9.3005
R1973 dvss.n326 dvss.n325 9.3005
R1974 dvss.n326 dvss.n147 9.3005
R1975 dvss.n332 dvss.n140 9.3005
R1976 dvss.n333 dvss.n332 9.3005
R1977 dvss.n332 dvss.n329 9.3005
R1978 dvss.n347 dvss.n346 9.3005
R1979 dvss.n346 dvss.n138 9.3005
R1980 dvss.n346 dvss.n345 9.3005
R1981 dvss.n560 dvss.n559 9.3005
R1982 dvss.n577 dvss.n576 9.3005
R1983 dvss.n576 dvss.n575 9.3005
R1984 dvss.n576 dvss.n125 9.3005
R1985 dvss.n582 dvss.n118 9.3005
R1986 dvss.n583 dvss.n582 9.3005
R1987 dvss.n582 dvss.n579 9.3005
R1988 dvss.n597 dvss.n596 9.3005
R1989 dvss.n596 dvss.n595 9.3005
R1990 dvss.n300 dvss.n299 9.3005
R1991 dvss.n156 dvss.n155 9.3005
R1992 dvss.n308 dvss.n307 9.3005
R1993 dvss.n153 dvss.n152 9.3005
R1994 dvss.n314 dvss.n313 9.3005
R1995 dvss.n312 dvss.n148 9.3005
R1996 dvss.n324 dvss.n323 9.3005
R1997 dvss.n322 dvss.n145 9.3005
R1998 dvss.n328 dvss.n144 9.3005
R1999 dvss.n335 dvss.n334 9.3005
R2000 dvss.n330 dvss.n141 9.3005
R2001 dvss.n343 dvss.n342 9.3005
R2002 dvss.n344 dvss.n137 9.3005
R2003 dvss.n349 dvss.n348 9.3005
R2004 dvss.n134 dvss.n133 9.3005
R2005 dvss.n558 dvss.n557 9.3005
R2006 dvss.n131 dvss.n130 9.3005
R2007 dvss.n564 dvss.n563 9.3005
R2008 dvss.n562 dvss.n126 9.3005
R2009 dvss.n574 dvss.n573 9.3005
R2010 dvss.n572 dvss.n123 9.3005
R2011 dvss.n578 dvss.n122 9.3005
R2012 dvss.n585 dvss.n584 9.3005
R2013 dvss.n580 dvss.n119 9.3005
R2014 dvss.n593 dvss.n592 9.3005
R2015 dvss.n594 dvss.n117 9.3005
R2016 dvss.n599 dvss.n598 9.3005
R2017 dvss.n654 dvss.n641 9.3005
R2018 dvss.n710 dvss.n709 9.3005
R2019 dvss.n708 dvss.n613 9.3005
R2020 dvss.n707 dvss.n706 9.3005
R2021 dvss.n705 dvss.n614 9.3005
R2022 dvss.n704 dvss.n703 9.3005
R2023 dvss.n702 dvss.n615 9.3005
R2024 dvss.n701 dvss.n700 9.3005
R2025 dvss.n699 dvss.n617 9.3005
R2026 dvss.n698 dvss.n697 9.3005
R2027 dvss.n696 dvss.n618 9.3005
R2028 dvss.n695 dvss.n694 9.3005
R2029 dvss.n693 dvss.n619 9.3005
R2030 dvss.n692 dvss.n691 9.3005
R2031 dvss.n688 dvss.n620 9.3005
R2032 dvss.n687 dvss.n686 9.3005
R2033 dvss.n685 dvss.n621 9.3005
R2034 dvss.n684 dvss.n683 9.3005
R2035 dvss.n682 dvss.n622 9.3005
R2036 dvss.n681 dvss.n680 9.3005
R2037 dvss.n679 dvss.n624 9.3005
R2038 dvss.n678 dvss.n677 9.3005
R2039 dvss.n676 dvss.n625 9.3005
R2040 dvss.n675 dvss.n674 9.3005
R2041 dvss.n673 dvss.n626 9.3005
R2042 dvss.n672 dvss.n671 9.3005
R2043 dvss.n670 dvss.n627 9.3005
R2044 dvss.n669 dvss.n629 9.3005
R2045 dvss.n668 dvss.n667 9.3005
R2046 dvss.n666 dvss.n631 9.3005
R2047 dvss.n665 dvss.n664 9.3005
R2048 dvss.n663 dvss.n632 9.3005
R2049 dvss.n662 dvss.n661 9.3005
R2050 dvss.n660 dvss.n635 9.3005
R2051 dvss.n659 dvss.n658 9.3005
R2052 dvss.n657 dvss.n636 9.3005
R2053 dvss.n656 dvss.n655 9.3005
R2054 dvss.n396 dvss.t13 9.18383
R2055 dvss.n396 dvss.t11 9.18383
R2056 dvss.n105 dvss.t53 9.18383
R2057 dvss.n105 dvss.t51 9.18383
R2058 dvss.n530 dvss.n517 8.79354
R2059 dvss.n993 dvss.n992 8.58924
R2060 dvss.t243 dvss.t210 8.43366
R2061 dvss.n80 dvss.t423 8.2655
R2062 dvss.n80 dvss.t380 8.2655
R2063 dvss.n79 dvss.t89 8.2655
R2064 dvss.n79 dvss.t425 8.2655
R2065 dvss.n776 dvss.t172 8.2655
R2066 dvss.n776 dvss.t225 8.2655
R2067 dvss.n777 dvss.t229 8.2655
R2068 dvss.n777 dvss.t116 8.2655
R2069 dvss.n778 dvss.t20 8.2655
R2070 dvss.n778 dvss.t184 8.2655
R2071 dvss.n749 dvss.n50 8.19036
R2072 dvss.n752 dvss.n93 8.18274
R2073 dvss.t407 dvss.t365 8.18274
R2074 dvss.n756 dvss.n738 8.18274
R2075 dvss.n1140 dvss.n796 8.15928
R2076 dvss.n1142 dvss.n1141 8.11042
R2077 dvss.n993 dvss.n961 8.03513
R2078 dvss.n1171 dvss.n1169 7.82362
R2079 dvss.n1433 dvss.n5 7.6805
R2080 dvss.n1167 dvss.n1166 7.13465
R2081 dvss.n1166 dvss.n1165 7.13465
R2082 dvss.n1164 dvss.n1163 7.13465
R2083 dvss.n1165 dvss.n1164 7.13465
R2084 dvss.n1158 dvss.n784 7.13465
R2085 dvss.n1162 dvss.n784 7.13465
R2086 dvss.n1161 dvss.n1160 7.13465
R2087 dvss.n1162 dvss.n1161 7.13465
R2088 dvss.n992 dvss.n991 7.01267
R2089 dvss.n1355 dvss.n1354 6.77697
R2090 dvss.n1071 dvss.n856 6.69588
R2091 dvss.n960 dvss.n954 6.4005
R2092 dvss.n1267 dvss.n1262 6.28553
R2093 dvss.n1433 dvss.n1432 6.26809
R2094 dvss.n531 dvss.n530 5.89963
R2095 dvss.n1131 dvss.n812 5.6454
R2096 dvss.n1072 dvss.n1071 5.61281
R2097 dvss.n454 dvss.n453 5.6005
R2098 dvss.n1273 dvss.n1272 5.51906
R2099 dvss.n466 dvss.n465 5.4005
R2100 dvss.n1258 dvss.n1256 5.13208
R2101 dvss.n1276 dvss.n1258 5.13208
R2102 dvss.n950 dvss.n815 5.12331
R2103 dvss.n546 dvss.n357 5.09503
R2104 dvss.n811 dvss.n795 5.08147
R2105 dvss.n764 dvss.n87 5.06981
R2106 dvss.n984 dvss.n983 5.05494
R2107 dvss.n1042 dvss.n903 5.02119
R2108 dvss.n764 dvss.n763 4.94307
R2109 dvss.n811 dvss.n810 4.86695
R2110 dvss.n1095 dvss.n1094 4.66041
R2111 dvss.n1270 dvss.n1269 4.65428
R2112 dvss.n173 dvss.n172 4.64132
R2113 dvss.n217 dvss.n216 4.64132
R2114 dvss.n311 dvss.n310 4.64111
R2115 dvss.n561 dvss.n560 4.64111
R2116 dvss.n1365 dvss.n30 4.6359
R2117 dvss.n1354 dvss.n1353 4.51815
R2118 dvss.n983 dvss.n934 4.46947
R2119 dvss.n1043 dvss.n1042 4.46947
R2120 dvss.n453 dvss.n452 4.38075
R2121 dvss.n492 dvss.n466 4.37879
R2122 dvss.n873 dvss.n864 4.36769
R2123 dvss.n934 dvss.n925 4.30062
R2124 dvss.n1252 dvss.n1250 4.29698
R2125 dvss.n1268 dvss.n1266 4.21607
R2126 dvss.n1266 dvss.n1265 4.14944
R2127 dvss.n1265 dvss.n1264 4.14944
R2128 dvss.t201 dvss.t350 4.09339
R2129 dvss.n1257 dvss.n1255 4.09141
R2130 dvss.n1259 dvss.n1257 4.09141
R2131 dvss.n726 dvss.n725 3.91448
R2132 dvss.n1294 dvss.n55 3.91161
R2133 dvss.n1055 dvss.n889 3.67161
R2134 dvss.n1022 dvss.n1019 3.66244
R2135 dvss.n1056 dvss.n1055 3.54509
R2136 dvss.n874 dvss.n873 3.50683
R2137 dvss.n1263 dvss.n1255 3.34378
R2138 dvss.n652 dvss.n651 3.27492
R2139 dvss.n990 dvss.n935 3.22833
R2140 dvss.n1045 dvss.n900 3.05772
R2141 dvss.n1044 dvss.n1043 3.05584
R2142 dvss.n1057 dvss.n888 2.94732
R2143 dvss.n532 dvss.n531 2.89441
R2144 dvss.n1130 dvss.n813 2.87229
R2145 dvss.n1073 dvss.n1072 2.86873
R2146 dvss.n1066 dvss.n1065 2.80414
R2147 dvss.n986 dvss.n985 2.61868
R2148 dvss.n989 dvss.n962 2.47323
R2149 dvss.n992 dvss.n989 2.47323
R2150 dvss.n1131 dvss.n1130 2.44756
R2151 dvss.n1169 dvss.n779 2.37019
R2152 dvss.n433 dvss.n399 2.35044
R2153 dvss.n440 dvss.n434 2.33839
R2154 dvss.n714 dvss.n713 2.19136
R2155 dvss.n418 dvss.n398 2.17408
R2156 dvss.n432 dvss.n431 2.09886
R2157 dvss.n879 dvss.n877 2.05207
R2158 dvss.n1021 dvss.n888 1.93399
R2159 dvss.n1120 dvss.n822 1.89703
R2160 dvss.n690 dvss.n688 1.86717
R2161 dvss.n1119 dvss.n1118 1.8605
R2162 dvss.n653 dvss.n652 1.8605
R2163 dvss.n1126 dvss.n1125 1.85699
R2164 dvss.n1220 dvss.t358 1.73948
R2165 dvss.n1210 dvss.t330 1.73948
R2166 dvss.n1190 dvss.t415 1.73948
R2167 dvss.n1240 dvss.t363 1.73948
R2168 dvss.n1057 dvss.n1056 1.72169
R2169 dvss.n1221 dvss.n1220 1.62652
R2170 dvss.n1222 dvss.n1221 1.62652
R2171 dvss.n1223 dvss.n1222 1.62652
R2172 dvss.n1224 dvss.n1223 1.62652
R2173 dvss.n1225 dvss.n1224 1.62652
R2174 dvss.n1226 dvss.n1225 1.62652
R2175 dvss.n1227 dvss.n1226 1.62652
R2176 dvss.n1228 dvss.n1227 1.62652
R2177 dvss.n1211 dvss.n1210 1.62652
R2178 dvss.n1212 dvss.n1211 1.62652
R2179 dvss.n1213 dvss.n1212 1.62652
R2180 dvss.n1214 dvss.n1213 1.62652
R2181 dvss.n1215 dvss.n1214 1.62652
R2182 dvss.n1216 dvss.n1215 1.62652
R2183 dvss.n1217 dvss.n1216 1.62652
R2184 dvss.n1218 dvss.n1217 1.62652
R2185 dvss.n1191 dvss.n1190 1.62652
R2186 dvss.n1192 dvss.n1191 1.62652
R2187 dvss.n1193 dvss.n1192 1.62652
R2188 dvss.n1194 dvss.n1193 1.62652
R2189 dvss.n1195 dvss.n1194 1.62652
R2190 dvss.n1196 dvss.n1195 1.62652
R2191 dvss.n1197 dvss.n1196 1.62652
R2192 dvss.n1198 dvss.n1197 1.62652
R2193 dvss.n1241 dvss.n1240 1.62652
R2194 dvss.n1242 dvss.n1241 1.62652
R2195 dvss.n1243 dvss.n1242 1.62652
R2196 dvss.n1244 dvss.n1243 1.62652
R2197 dvss.n1245 dvss.n1244 1.62652
R2198 dvss.n1246 dvss.n1245 1.62652
R2199 dvss.n1247 dvss.n1246 1.62652
R2200 dvss.n1248 dvss.n1247 1.62652
R2201 dvss.n1274 dvss.n1273 1.56886
R2202 dvss.n1275 dvss.n1274 1.56886
R2203 dvss.n1100 dvss.n1099 1.5505
R2204 dvss.n1252 dvss.n1251 1.50955
R2205 dvss.n1069 dvss.n1068 1.49704
R2206 dvss.n1117 avss 1.48104
R2207 dvss.n711 dvss.n710 1.45077
R2208 dvss.n411 dvss.n399 1.44956
R2209 dvss.n611 dvss 1.44157
R2210 dvss.n859 dvss.n842 1.32133
R2211 dvss.n861 dvss.n823 1.31102
R2212 dvss.n1434 dvss.n4 1.30418
R2213 dvss.n612 dvss.n611 1.29478
R2214 dvss.n724 dvss.n723 1.24591
R2215 dvss.n1097 avss 1.23982
R2216 dvss.n434 dvss.n398 1.23022
R2217 dvss.n434 dvss.n433 1.22373
R2218 dvss.n723 dvss.n722 1.22095
R2219 dvss.n1280 dvss.n1279 1.20521
R2220 dvss.n1116 dvss.n1115 1.19172
R2221 dvss.n1219 dvss.n1218 1.16356
R2222 dvss.n1199 dvss.n1198 1.16356
R2223 dvss.n1249 dvss.n1248 1.16047
R2224 dvss.n1229 dvss.n1228 1.1604
R2225 dvss.n1279 dvss.n1278 1.13422
R2226 dvss.n1278 dvss.n1277 1.13422
R2227 dvss.n1289 dvss.n1288 1.09721
R2228 dvss.n1045 dvss.n1044 1.09236
R2229 dvss.n1069 dvss.n848 1.06941
R2230 dvss.n653 dvss.n4 1.0534
R2231 dvss.n531 dvss.n108 1.01717
R2232 dvss.n1154 dvss.n1153 0.969941
R2233 dvss.n1067 dvss.n1066 0.957122
R2234 dvss.n1018 dvss.n1017 0.893523
R2235 dvss.n867 dvss.n863 0.845955
R2236 dvss.n1096 dvss.n1095 0.845955
R2237 dvss.n901 dvss.n890 0.841376
R2238 dvss.n1283 dvss.n1252 0.808157
R2239 dvss.n653 dvss.n642 0.776443
R2240 dvss.n1361 dvss.n1359 0.753441
R2241 dvss dvss.n4 0.733375
R2242 dvss.n1101 dvss.n840 0.731929
R2243 dvss.n1157 dvss.n1156 0.714663
R2244 dvss.n611 dvss 0.71054
R2245 dvss.n1096 dvss.n842 0.686469
R2246 dvss.n1285 dvss.t319 0.685626
R2247 dvss.n1288 dvss 0.679512
R2248 dvss.n1024 dvss.n1023 0.672416
R2249 dvss.n1286 dvss.t207 0.659973
R2250 dvss.n1075 dvss.n1074 0.650441
R2251 dvss.n1129 dvss.n815 0.649705
R2252 dvss.n773 dvss.n772 0.647619
R2253 dvss.n1288 dvss.n1287 0.626581
R2254 dvss.n785 dvss.n26 0.620568
R2255 dvss.t248 dvss.t245 0.620568
R2256 dvss.t239 dvss.t157 0.620568
R2257 dvss.t238 dvss.t124 0.620568
R2258 dvss.t140 dvss.t9 0.620568
R2259 dvss.t242 dvss.t342 0.620568
R2260 dvss.t179 dvss.t367 0.620568
R2261 dvss.t72 dvss.t29 0.620568
R2262 dvss.t34 dvss.t106 0.620568
R2263 dvss.t27 dvss.t414 0.620568
R2264 dvss.t38 dvss.t62 0.620568
R2265 dvss.t432 dvss.t400 0.620568
R2266 dvss.t118 dvss.t338 0.620568
R2267 dvss.n1165 dvss.n1162 0.620568
R2268 dvss.t437 dvss.t39 0.620568
R2269 dvss.t178 dvss.t174 0.620568
R2270 dvss.t177 dvss.t279 0.620568
R2271 dvss.t85 dvss.t339 0.620568
R2272 dvss.t249 dvss.t397 0.620568
R2273 dvss.t262 dvss.t315 0.620568
R2274 dvss.t247 dvss.t316 0.620568
R2275 dvss.t28 dvss.t123 0.620568
R2276 dvss.t383 dvss.t409 0.620568
R2277 dvss.t436 dvss.t173 0.620568
R2278 dvss.t435 dvss.t4 0.620568
R2279 dvss.t63 dvss.t117 0.620568
R2280 dvss.n1147 dvss.n787 0.620568
R2281 dvss.n1093 dvss.n842 0.6205
R2282 dvss.n1154 dvss.n779 0.617214
R2283 dvss.n1068 dvss.n863 0.606103
R2284 dvss.n1098 dvss.n1097 0.604749
R2285 dvss.n770 dvss.n769 0.603757
R2286 dvss.n357 dvss.n104 0.603227
R2287 dvss.n1074 dvss.n1070 0.593683
R2288 dvss.n1284 dvss.n1171 0.584781
R2289 dvss.n815 dvss.n813 0.584691
R2290 dvss.n1115 dvss.n1114 0.582318
R2291 dvss.n771 dvss.n770 0.573586
R2292 dvss.n861 avss 0.566822
R2293 dvss.n1284 dvss.n1283 0.53923
R2294 dvss.n859 dvss.n858 0.517167
R2295 dvss.n1229 dvss.n1219 0.501662
R2296 dvss.n1170 dvss.t474 0.487968
R2297 dvss.n1008 dvss.n935 0.457643
R2298 dvss.n1171 dvss.n1170 0.448591
R2299 dvss.n1169 dvss.n1168 0.407877
R2300 dvss.n1099 dvss.n1098 0.406136
R2301 dvss.n714 dvss.n103 0.404873
R2302 dvss.n433 dvss.n432 0.404848
R2303 dvss.n1116 dvss.n824 0.398755
R2304 dvss.n860 dvss.n859 0.39776
R2305 dvss.n770 dvss.n81 0.396762
R2306 dvss.n1067 dvss.n864 0.389389
R2307 dvss.n860 dvss.n824 0.388725
R2308 dvss.n775 dvss.n774 0.38836
R2309 dvss.n1019 dvss.n925 0.386852
R2310 dvss.n1285 dvss.t467 0.372324
R2311 dvss.n1286 dvss.t480 0.368665
R2312 dvss.n1022 dvss.n1021 0.358192
R2313 dvss dvss.n653 0.356294
R2314 dvss.n1023 dvss.n900 0.353256
R2315 dvss.n1270 dvss.n1262 0.344944
R2316 dvss.n1129 dvss.n1128 0.335899
R2317 dvss.n1118 dvss.n1117 0.32778
R2318 dvss.n1118 dvss.n822 0.323689
R2319 dvss.n1251 dvss.t479 0.315839
R2320 dvss.n1020 dvss.n900 0.3105
R2321 dvss.n1287 dvss.n1285 0.310127
R2322 dvss.n716 dvss.n715 0.30764
R2323 dvss.n1153 dvss.n1152 0.307378
R2324 dvss.n1098 dvss.n840 0.3005
R2325 dvss.n1434 dvss.n1433 0.3005
R2326 dvss.n981 dvss.n888 0.298417
R2327 dvss.n812 dvss.n811 0.293439
R2328 dvss.n1294 dvss.n1293 0.284911
R2329 dvss.n862 dvss.n860 0.28415
R2330 dvss.n1156 dvss.n1155 0.275178
R2331 dvss.n1058 dvss.n1057 0.266214
R2332 avss dvss.n1116 0.260623
R2333 dvss.n864 dvss.n863 0.256966
R2334 dvss.n742 dvss.n88 0.253965
R2335 dvss.n744 dvss.n743 0.253965
R2336 dvss.n772 dvss.n771 0.240989
R2337 dvss.n377 dvss.n370 0.238561
R2338 dvss.n493 dvss.n462 0.238561
R2339 dvss.n1249 dvss.n1239 0.236669
R2340 dvss.n1199 dvss.n1189 0.23559
R2341 dvss.n774 dvss.n773 0.227866
R2342 dvss.n719 dvss.n718 0.227486
R2343 dvss.n1291 dvss.n1290 0.226323
R2344 dvss.n1155 dvss.n1154 0.221929
R2345 dvss.n1292 dvss.n1291 0.221179
R2346 dvss.n1290 dvss.n1289 0.220665
R2347 dvss.n2 dvss.n1 0.214786
R2348 dvss.n1250 dvss.n1249 0.214159
R2349 dvss.n720 dvss.n81 0.213219
R2350 dvss.n722 dvss.n716 0.210077
R2351 dvss.n1056 dvss.n886 0.207167
R2352 dvss.n1209 dvss.n1199 0.203775
R2353 dvss.n1097 dvss.n1096 0.20273
R2354 dvss.n1152 dvss.n3 0.20222
R2355 dvss.n1251 dvss.t170 0.201112
R2356 dvss.n441 dvss.n440 0.195503
R2357 dvss.n1127 dvss.n1126 0.179346
R2358 dvss.n720 dvss.n719 0.178167
R2359 dvss.n1230 dvss.n1229 0.177752
R2360 avss dvss.n1069 0.173899
R2361 dvss.n1287 dvss.n1286 0.171
R2362 dvss.n612 dvss.n108 0.170624
R2363 dvss.n107 dvss.n106 0.165438
R2364 dvss.n1059 dvss.n886 0.163557
R2365 dvss.n715 dvss.n714 0.16209
R2366 dvss.n1219 dvss.n1209 0.15883
R2367 dvss.n385 dvss.n384 0.157363
R2368 dvss.n386 dvss.n385 0.157363
R2369 dvss.n387 dvss.n386 0.157363
R2370 dvss.n388 dvss.n387 0.157363
R2371 dvss.n389 dvss.n388 0.157363
R2372 dvss.n450 dvss.n449 0.157363
R2373 dvss.n449 dvss.n448 0.157363
R2374 dvss.n448 dvss.n447 0.157363
R2375 dvss.n447 dvss.n446 0.157363
R2376 dvss.n446 dvss.n445 0.157363
R2377 dvss.n474 dvss.n473 0.157363
R2378 dvss.n475 dvss.n474 0.157363
R2379 dvss.n476 dvss.n475 0.157363
R2380 dvss.n477 dvss.n476 0.157363
R2381 dvss.n478 dvss.n477 0.157363
R2382 dvss.n490 dvss.n489 0.157363
R2383 dvss.n489 dvss.n488 0.157363
R2384 dvss.n488 dvss.n487 0.157363
R2385 dvss.n487 dvss.n486 0.157363
R2386 dvss.n486 dvss.n485 0.157363
R2387 dvss.n485 dvss.n103 0.157363
R2388 dvss.n1117 dvss.n823 0.152695
R2389 dvss.n1128 dvss.n812 0.148401
R2390 dvss.n1435 dvss.n1434 0.129071
R2391 dvss.n444 dvss.n442 0.122553
R2392 dvss.n711 dvss.n612 0.119023
R2393 dvss dvss.n1284 0.118752
R2394 dvss.n451 dvss.n389 0.115696
R2395 dvss.n491 dvss.n478 0.115696
R2396 dvss.n1228 dvss.t348 0.113463
R2397 dvss.n1227 dvss.t347 0.113463
R2398 dvss.n1226 dvss.t362 0.113463
R2399 dvss.n1225 dvss.t361 0.113463
R2400 dvss.n1224 dvss.t352 0.113463
R2401 dvss.n1223 dvss.t343 0.113463
R2402 dvss.n1222 dvss.t355 0.113463
R2403 dvss.n1221 dvss.t364 0.113463
R2404 dvss.n1220 dvss.t344 0.113463
R2405 dvss.n1218 dvss.t194 0.113463
R2406 dvss.n1217 dvss.t193 0.113463
R2407 dvss.n1216 dvss.t197 0.113463
R2408 dvss.n1215 dvss.t196 0.113463
R2409 dvss.n1214 dvss.t195 0.113463
R2410 dvss.n1213 dvss.t198 0.113463
R2411 dvss.n1212 dvss.t333 0.113463
R2412 dvss.n1211 dvss.t331 0.113463
R2413 dvss.n1210 dvss.t332 0.113463
R2414 dvss.n1198 dvss.t325 0.113463
R2415 dvss.n1197 dvss.t324 0.113463
R2416 dvss.n1196 dvss.t328 0.113463
R2417 dvss.n1195 dvss.t327 0.113463
R2418 dvss.n1194 dvss.t326 0.113463
R2419 dvss.n1193 dvss.t329 0.113463
R2420 dvss.n1192 dvss.t418 0.113463
R2421 dvss.n1191 dvss.t416 0.113463
R2422 dvss.n1190 dvss.t417 0.113463
R2423 dvss.n1248 dvss.t357 0.113463
R2424 dvss.n1247 dvss.t356 0.113463
R2425 dvss.n1246 dvss.t346 0.113463
R2426 dvss.n1245 dvss.t345 0.113463
R2427 dvss.n1244 dvss.t359 0.113463
R2428 dvss.n1243 dvss.t353 0.113463
R2429 dvss.n1242 dvss.t360 0.113463
R2430 dvss.n1241 dvss.t349 0.113463
R2431 dvss.n1240 dvss.t354 0.113463
R2432 dvss.n106 dvss 0.112015
R2433 dvss.n1099 dvss.n824 0.109693
R2434 dvss.n712 dvss.n711 0.107057
R2435 dvss.n858 dvss.n844 0.106285
R2436 dvss.n1435 dvss.n3 0.105659
R2437 dvss.n452 dvss.n451 0.105151
R2438 dvss.n492 dvss.n491 0.105151
R2439 dvss.n1172 dvss.t447 0.10275
R2440 dvss.n1181 dvss.t482 0.10275
R2441 dvss.n1200 dvss.t472 0.10275
R2442 dvss.n1231 dvss.t455 0.10275
R2443 dvss.n445 dvss.n444 0.102624
R2444 dvss.n439 dvss.n438 0.100225
R2445 dvss dvss.n1435 0.0930926
R2446 dvss.n1365 dvss.n1364 0.0918107
R2447 dvss.n642 dvss 0.0911863
R2448 dvss.n1256 dvss.n1254 0.0907913
R2449 dvss.n1070 avss 0.0896768
R2450 dvss.n1055 dvss.n1054 0.0866111
R2451 dvss dvss.n81 0.084875
R2452 dvss.n1209 dvss.n1208 0.0788906
R2453 dvss.n713 dvss.n104 0.0765474
R2454 dvss.n1128 dvss.n1127 0.0758817
R2455 dvss.n1293 dvss.n775 0.0756029
R2456 dvss.n715 dvss 0.0731595
R2457 dvss.n442 dvss.n441 0.0723713
R2458 dvss.n1269 dvss.n1268 0.0709545
R2459 dvss.n1263 dvss.n1253 0.0704248
R2460 dvss.n1170 dvss.t396 0.069705
R2461 dvss.n1173 dvss.n1172 0.06865
R2462 dvss.n1174 dvss.n1173 0.06865
R2463 dvss.n1175 dvss.n1174 0.06865
R2464 dvss.n1176 dvss.n1175 0.06865
R2465 dvss.n1177 dvss.n1176 0.06865
R2466 dvss.n1178 dvss.n1177 0.06865
R2467 dvss.n1179 dvss.n1178 0.06865
R2468 dvss.n1180 dvss.n1179 0.06865
R2469 dvss.n1182 dvss.n1181 0.06865
R2470 dvss.n1183 dvss.n1182 0.06865
R2471 dvss.n1184 dvss.n1183 0.06865
R2472 dvss.n1185 dvss.n1184 0.06865
R2473 dvss.n1186 dvss.n1185 0.06865
R2474 dvss.n1187 dvss.n1186 0.06865
R2475 dvss.n1188 dvss.n1187 0.06865
R2476 dvss.n1189 dvss.n1188 0.06865
R2477 dvss.n1201 dvss.n1200 0.06865
R2478 dvss.n1202 dvss.n1201 0.06865
R2479 dvss.n1203 dvss.n1202 0.06865
R2480 dvss.n1204 dvss.n1203 0.06865
R2481 dvss.n1205 dvss.n1204 0.06865
R2482 dvss.n1206 dvss.n1205 0.06865
R2483 dvss.n1207 dvss.n1206 0.06865
R2484 dvss.n1208 dvss.n1207 0.06865
R2485 dvss.n1232 dvss.n1231 0.06865
R2486 dvss.n1233 dvss.n1232 0.06865
R2487 dvss.n1234 dvss.n1233 0.06865
R2488 dvss.n1235 dvss.n1234 0.06865
R2489 dvss.n1236 dvss.n1235 0.06865
R2490 dvss.n1237 dvss.n1236 0.06865
R2491 dvss.n1238 dvss.n1237 0.06865
R2492 dvss.n1239 dvss.n1238 0.06865
R2493 dvss.n442 dvss.n397 0.0660593
R2494 dvss.n1230 dvss.n1180 0.0632125
R2495 dvss dvss.n1365 0.0615076
R2496 dvss.n1318 dvss.n1317 0.0611061
R2497 dvss.n1319 dvss.n1318 0.0611061
R2498 dvss.n1319 dvss.n44 0.0611061
R2499 dvss.n1323 dvss.n44 0.0611061
R2500 dvss.n1324 dvss.n1323 0.0611061
R2501 dvss.n1325 dvss.n1324 0.0611061
R2502 dvss.n1325 dvss.n41 0.0611061
R2503 dvss.n1329 dvss.n41 0.0611061
R2504 dvss.n1330 dvss.n1329 0.0611061
R2505 dvss.n1331 dvss.n1330 0.0611061
R2506 dvss.n1331 dvss.n39 0.0611061
R2507 dvss.n1336 dvss.n39 0.0611061
R2508 dvss.n1337 dvss.n1336 0.0611061
R2509 dvss.n1338 dvss.n1337 0.0611061
R2510 dvss.n1338 dvss.n37 0.0611061
R2511 dvss.n1342 dvss.n37 0.0611061
R2512 dvss.n1343 dvss.n1342 0.0611061
R2513 dvss.n1344 dvss.n1343 0.0611061
R2514 dvss.n1344 dvss.n35 0.0611061
R2515 dvss.n1349 dvss.n35 0.0611061
R2516 dvss.n1350 dvss.n1349 0.0611061
R2517 dvss.n1351 dvss.n1350 0.0611061
R2518 dvss.n1356 dvss.n33 0.0611061
R2519 dvss.n1357 dvss.n1356 0.0611061
R2520 dvss.n1358 dvss.n1357 0.0611061
R2521 dvss.n1358 dvss.n31 0.0611061
R2522 dvss.n1364 dvss.n31 0.0611061
R2523 dvss.n1373 dvss.n1367 0.0611061
R2524 dvss.n1373 dvss.n1372 0.0611061
R2525 dvss.n706 dvss.n613 0.0550455
R2526 dvss.n706 dvss.n705 0.0550455
R2527 dvss.n705 dvss.n704 0.0550455
R2528 dvss.n704 dvss.n615 0.0550455
R2529 dvss.n700 dvss.n615 0.0550455
R2530 dvss.n700 dvss.n699 0.0550455
R2531 dvss.n699 dvss.n698 0.0550455
R2532 dvss.n698 dvss.n618 0.0550455
R2533 dvss.n694 dvss.n618 0.0550455
R2534 dvss.n694 dvss.n693 0.0550455
R2535 dvss.n693 dvss.n692 0.0550455
R2536 dvss.n692 dvss.n620 0.0550455
R2537 dvss.n686 dvss.n620 0.0550455
R2538 dvss.n686 dvss.n685 0.0550455
R2539 dvss.n685 dvss.n684 0.0550455
R2540 dvss.n684 dvss.n622 0.0550455
R2541 dvss.n680 dvss.n622 0.0550455
R2542 dvss.n680 dvss.n679 0.0550455
R2543 dvss.n679 dvss.n678 0.0550455
R2544 dvss.n678 dvss.n625 0.0550455
R2545 dvss.n674 dvss.n625 0.0550455
R2546 dvss.n674 dvss.n673 0.0550455
R2547 dvss.n672 dvss.n627 0.0550455
R2548 dvss.n629 dvss.n627 0.0550455
R2549 dvss.n667 dvss.n629 0.0550455
R2550 dvss.n667 dvss.n666 0.0550455
R2551 dvss.n666 dvss.n665 0.0550455
R2552 dvss.n665 dvss.n632 0.0550455
R2553 dvss.n661 dvss.n632 0.0550455
R2554 dvss.n661 dvss.n660 0.0550455
R2555 dvss.n660 dvss.n659 0.0550455
R2556 dvss.n659 dvss.n636 0.0550455
R2557 dvss.n655 dvss.n636 0.0550455
R2558 dvss.n718 dvss.n717 0.054997
R2559 dvss.n308 dvss.n155 0.0533634
R2560 dvss.n313 dvss.n312 0.0533634
R2561 dvss.n344 dvss.n343 0.0533634
R2562 dvss.n558 dvss.n133 0.0533634
R2563 dvss.n563 dvss.n562 0.0533634
R2564 dvss.n594 dvss.n593 0.0533634
R2565 dvss.n721 dvss.n720 0.0533607
R2566 dvss.n169 dvss.n164 0.0522241
R2567 dvss.n175 dvss.n174 0.0522241
R2568 dvss.n201 dvss.n200 0.0522241
R2569 dvss.n212 dvss.n211 0.0522241
R2570 dvss.n226 dvss.n218 0.0522241
R2571 dvss.n607 dvss.n110 0.0522241
R2572 dvss.n440 dvss.n439 0.0510502
R2573 dvss.n1371 dvss 0.0503737
R2574 dvss.n1020 avss 0.0500072
R2575 dvss.n329 dvss.n328 0.0484075
R2576 dvss.n579 dvss.n578 0.0484075
R2577 dvss.n1293 dvss.n1292 0.0483395
R2578 dvss.n195 dvss.n187 0.047375
R2579 dvss.n237 dvss.n232 0.047375
R2580 dvss.n328 dvss.n327 0.0451035
R2581 dvss.n578 dvss.n577 0.0451035
R2582 dvss.n187 dvss.n186 0.0441422
R2583 dvss.n232 dvss.n231 0.0441422
R2584 dvss.n713 dvss.n712 0.0428497
R2585 dvss.n451 dvss.n450 0.0421667
R2586 dvss.n491 dvss.n490 0.0421667
R2587 dvss.n862 dvss.n861 0.0421667
R2588 dvss.n1372 dvss.n1371 0.0415354
R2589 dvss.n1283 dvss.n1282 0.0392931
R2590 dvss.n312 dvss.n147 0.0351916
R2591 dvss.n334 dvss.n333 0.0351916
R2592 dvss.n348 dvss.n347 0.0351916
R2593 dvss.n562 dvss.n125 0.0351916
R2594 dvss.n584 dvss.n583 0.0351916
R2595 dvss.n1172 dvss.t448 0.0346
R2596 dvss.n1173 dvss.t478 0.0346
R2597 dvss.n1174 dvss.t462 0.0346
R2598 dvss.n1175 dvss.t463 0.0346
R2599 dvss.n1176 dvss.t449 0.0346
R2600 dvss.n1177 dvss.t450 0.0346
R2601 dvss.n1178 dvss.t475 0.0346
R2602 dvss.n1179 dvss.t458 0.0346
R2603 dvss.n1180 dvss.t459 0.0346
R2604 dvss.n1181 dvss.t483 0.0346
R2605 dvss.n1182 dvss.t471 0.0346
R2606 dvss.n1183 dvss.t453 0.0346
R2607 dvss.n1184 dvss.t454 0.0346
R2608 dvss.n1185 dvss.t442 0.0346
R2609 dvss.n1186 dvss.t444 0.0346
R2610 dvss.n1187 dvss.t468 0.0346
R2611 dvss.n1188 dvss.t451 0.0346
R2612 dvss.n1189 dvss.t452 0.0346
R2613 dvss.n1200 dvss.t473 0.0346
R2614 dvss.n1201 dvss.t464 0.0346
R2615 dvss.n1202 dvss.t443 0.0346
R2616 dvss.n1203 dvss.t445 0.0346
R2617 dvss.n1204 dvss.t476 0.0346
R2618 dvss.n1205 dvss.t477 0.0346
R2619 dvss.n1206 dvss.t457 0.0346
R2620 dvss.n1207 dvss.t484 0.0346
R2621 dvss.n1208 dvss.t440 0.0346
R2622 dvss.n1231 dvss.t456 0.0346
R2623 dvss.n1232 dvss.t446 0.0346
R2624 dvss.n1233 dvss.t469 0.0346
R2625 dvss.n1234 dvss.t470 0.0346
R2626 dvss.n1235 dvss.t460 0.0346
R2627 dvss.n1236 dvss.t461 0.0346
R2628 dvss.n1237 dvss.t441 0.0346
R2629 dvss.n1238 dvss.t465 0.0346
R2630 dvss.n1239 dvss.t466 0.0346
R2631 dvss.n181 dvss.n175 0.034444
R2632 dvss.n196 dvss.n188 0.034444
R2633 dvss.n210 dvss.n202 0.034444
R2634 dvss.n227 dvss.n226 0.034444
R2635 dvss.n236 dvss.n235 0.034444
R2636 dvss.n1024 dvss.n1022 0.0340958
R2637 dvss.n598 dvss.n595 0.0335396
R2638 dvss.n608 dvss.n109 0.0328276
R2639 dvss.n309 dvss.n153 0.0318877
R2640 dvss.n325 dvss.n145 0.0318877
R2641 dvss.n343 dvss.n140 0.0318877
R2642 dvss.n559 dvss.n131 0.0318877
R2643 dvss.n575 dvss.n123 0.0318877
R2644 dvss.n593 dvss.n118 0.0318877
R2645 dvss.n170 dvss.n168 0.0312112
R2646 dvss.n183 dvss.n180 0.0312112
R2647 dvss.n200 dvss.n199 0.0312112
R2648 dvss.n214 dvss.n213 0.0312112
R2649 dvss.n228 dvss.n225 0.0312112
R2650 dvss.n240 dvss.n110 0.0312112
R2651 dvss.n1317 dvss 0.030803
R2652 dvss.n1351 dvss 0.030803
R2653 dvss dvss.n33 0.030803
R2654 dvss.n1366 dvss 0.030803
R2655 dvss dvss.n1366 0.030803
R2656 dvss.n1367 dvss 0.030803
R2657 dvss.n299 dvss.n298 0.0302357
R2658 dvss.n163 dvss.n161 0.0295948
R2659 dvss.n311 dvss.n153 0.0290415
R2660 dvss.n561 dvss.n131 0.0290415
R2661 dvss.n173 dvss.n168 0.0284381
R2662 dvss.n217 dvss.n213 0.0284381
R2663 dvss.n710 dvss 0.0277727
R2664 dvss.n613 dvss 0.0277727
R2665 dvss.n673 dvss 0.0277727
R2666 dvss dvss.n672 0.0277727
R2667 dvss.n655 dvss 0.0277727
R2668 dvss dvss.n654 0.0277727
R2669 dvss.n654 dvss 0.0277727
R2670 dvss.n1272 dvss.n1271 0.0266972
R2671 dvss.n313 dvss.n311 0.0257376
R2672 dvss.n563 dvss.n561 0.0257376
R2673 dvss.n174 dvss.n173 0.0252053
R2674 dvss.n218 dvss.n217 0.0252053
R2675 dvss.n1370 dvss 0.0246935
R2676 dvss.n298 dvss.n155 0.0236278
R2677 dvss.n164 dvss.n163 0.0231293
R2678 dvss.n309 dvss.n308 0.0219758
R2679 dvss.n325 dvss.n324 0.0219758
R2680 dvss.n330 dvss.n140 0.0219758
R2681 dvss dvss.n138 0.0219758
R2682 dvss.n559 dvss.n558 0.0219758
R2683 dvss.n575 dvss.n574 0.0219758
R2684 dvss.n580 dvss.n118 0.0219758
R2685 dvss.n170 dvss.n169 0.0215129
R2686 dvss.n183 dvss.n182 0.0215129
R2687 dvss.n199 dvss.n194 0.0215129
R2688 dvss.n207 dvss 0.0215129
R2689 dvss.n214 dvss.n212 0.0215129
R2690 dvss.n228 dvss.n224 0.0215129
R2691 dvss.n241 dvss.n240 0.0215129
R2692 dvss.n595 dvss.n594 0.0203238
R2693 dvss.n597 dvss 0.0203238
R2694 dvss.n608 dvss.n607 0.0198966
R2695 dvss dvss.n610 0.0198966
R2696 dvss.n1281 dvss.n1280 0.0196358
R2697 dvss.n324 dvss.n147 0.0186718
R2698 dvss.n333 dvss.n330 0.0186718
R2699 dvss.n345 dvss 0.0186718
R2700 dvss.n347 dvss.n133 0.0186718
R2701 dvss.n574 dvss.n125 0.0186718
R2702 dvss.n583 dvss.n580 0.0186718
R2703 dvss.n182 dvss.n181 0.0182802
R2704 dvss.n196 dvss.n194 0.0182802
R2705 dvss dvss.n206 0.0182802
R2706 dvss.n211 dvss.n210 0.0182802
R2707 dvss.n227 dvss.n224 0.0182802
R2708 dvss.n241 dvss.n235 0.0182802
R2709 dvss.n397 dvss.n104 0.0180319
R2710 dvss.n1070 dvss.n862 0.0176494
R2711 dvss.n1371 dvss.n1370 0.016125
R2712 dvss.n1021 dvss.n1020 0.0146129
R2713 dvss dvss.n2 0.0143889
R2714 dvss.n1127 avss 0.0133817
R2715 dvss.n108 dvss.n107 0.0129481
R2716 dvss.n452 dvss.n377 0.0125063
R2717 dvss.n493 dvss.n492 0.0125063
R2718 dvss.n823 avss 0.0119504
R2719 dvss.n299 dvss.n296 0.0104119
R2720 dvss.n161 dvss.n160 0.0101983
R2721 dvss.n1068 dvss.n1067 0.00875991
R2722 dvss.n327 dvss.n145 0.00875991
R2723 dvss.n345 dvss.n344 0.00875991
R2724 dvss.n577 dvss.n123 0.00875991
R2725 dvss.n186 dvss.n180 0.0085819
R2726 dvss.n206 dvss.n201 0.0085819
R2727 dvss.n231 dvss.n225 0.0085819
R2728 dvss.n598 dvss.n597 0.00710793
R2729 dvss.n610 dvss.n109 0.00696552
R2730 dvss.n722 dvss.n721 0.00671891
R2731 dvss.n1282 dvss.n1281 0.00626923
R2732 dvss.n334 dvss.n329 0.00545595
R2733 dvss.n348 dvss.n138 0.00545595
R2734 dvss.n584 dvss.n579 0.00545595
R2735 dvss.n195 dvss.n188 0.00534914
R2736 dvss.n207 dvss.n202 0.00534914
R2737 dvss.n237 dvss.n236 0.00534914
R2738 dvss.n1250 dvss.n1230 0.00291667
R2739 x2.VT2.t11 x2.VT2.n7 291.022
R2740 x2.VT2.n0 x2.VT2.t9 290.637
R2741 x2.VT2.n0 x2.VT2.t11 290.637
R2742 x2.VT2.t9 x2.VT2.n7 290.637
R2743 x2.VT2.n5 x2.VT2.t10 256.478
R2744 x2.VT2.t10 x2.VT2.n3 256.454
R2745 x2.VT2.n5 x2.VT2.t8 256.094
R2746 x2.VT2.t8 x2.VT2.n3 256.094
R2747 x2.VT2.n9 x2.VT2.n6 204.623
R2748 x2.VT2.n1 x2.VT2.n4 199.334
R2749 x2.VT2.n4 x2.VT2.t6 34.8005
R2750 x2.VT2.n4 x2.VT2.t4 34.8005
R2751 x2.VT2.n6 x2.VT2.t5 28.5655
R2752 x2.VT2.n6 x2.VT2.t7 28.5655
R2753 x2.VT2 x2.VT2.n1 5.87598
R2754 x2.VT2 x2.VT2.n9 1.25513
R2755 x2.VT2.n1 x2.VT2.n5 1.21382
R2756 x2.VT2.n9 x2.VT2.n8 0.799792
R2757 x2.VT2.t0 x2.VT2.n2 0.69766
R2758 x2.VT2.t1 x2.VT2.t3 0.489041
R2759 x2.VT2.n8 x2.VT2.n7 0.412638
R2760 x2.VT2.n0 x2.VT2.t2 16.4059
R2761 x2.VT2.n8 x2.VT2.n0 1.30841
R2762 x2.VT2.t2 x2.VT2.t1 0.672434
R2763 x2.VT2.t0 x2.VT2.t2 0.61243
R2764 x2.VT2.n1 x2.VT2.n3 0.513879
R2765 dvdd.n102 dvdd.n100 5954.12
R2766 dvdd.n103 dvdd.n100 5954.12
R2767 dvdd.n103 dvdd.n99 5954.12
R2768 dvdd.n102 dvdd.n99 5954.12
R2769 dvdd.n114 dvdd.n111 5954.12
R2770 dvdd.n114 dvdd.n112 5954.12
R2771 dvdd.n115 dvdd.n111 5954.12
R2772 dvdd.n115 dvdd.n112 5954.12
R2773 dvdd.n516 dvdd.n493 2258.82
R2774 dvdd.n516 dvdd.n494 2258.82
R2775 dvdd.n508 dvdd.n499 2258.82
R2776 dvdd.n594 dvdd.n589 2177.65
R2777 dvdd.n596 dvdd.n589 2177.65
R2778 dvdd.n453 dvdd.n449 2177.65
R2779 dvdd.n451 dvdd.n449 2177.65
R2780 dvdd.n603 dvdd.n602 1994.12
R2781 dvdd.n519 dvdd.n490 1994.12
R2782 dvdd.n520 dvdd.n519 1994.12
R2783 dvdd.n284 dvdd 1968.26
R2784 dvdd.n386 dvdd.n346 1838.82
R2785 dvdd.n549 dvdd.n312 1838.82
R2786 dvdd.n423 dvdd.n417 1838.82
R2787 dvdd.n423 dvdd.n415 1838.82
R2788 dvdd.n380 dvdd.n351 1697.65
R2789 dvdd.n377 dvdd.n356 1697.65
R2790 dvdd.n373 dvdd.n356 1697.65
R2791 dvdd.n506 dvdd.n505 1648.24
R2792 dvdd.n506 dvdd.n498 1648.24
R2793 dvdd.n153 dvdd.n150 1514.12
R2794 dvdd.n155 dvdd.n150 1514.12
R2795 dvdd.n161 dvdd.n147 1514.12
R2796 dvdd.n159 dvdd.n147 1514.12
R2797 dvdd.n274 dvdd.n269 1443.53
R2798 dvdd.n274 dvdd.n270 1443.53
R2799 dvdd.n272 dvdd.n269 1443.53
R2800 dvdd.n272 dvdd.n270 1443.53
R2801 dvdd.n591 dvdd.n583 1436.47
R2802 dvdd.n591 dvdd.n590 1436.47
R2803 dvdd.n609 dvdd.n584 1436.47
R2804 dvdd.n609 dvdd.n586 1436.47
R2805 dvdd.n524 dvdd.n461 1436.47
R2806 dvdd.n524 dvdd.n463 1436.47
R2807 dvdd.n458 dvdd.n447 1436.47
R2808 dvdd.n458 dvdd.n443 1436.47
R2809 dvdd.n455 dvdd.n446 1436.47
R2810 dvdd.n455 dvdd.n442 1436.47
R2811 dvdd.n507 dvdd.n494 1431.25
R2812 dvdd.n508 dvdd.n507 1431.25
R2813 dvdd.n373 dvdd.n368 1231.76
R2814 dvdd.n478 dvdd.n472 1110.52
R2815 dvdd.n478 dvdd.n473 1110.52
R2816 dvdd.n476 dvdd.n473 1110.52
R2817 dvdd.n476 dvdd.n472 1110.52
R2818 dvdd.n384 dvdd.n348 960
R2819 dvdd.n384 dvdd.n340 960
R2820 dvdd.n398 dvdd.n340 960
R2821 dvdd.n398 dvdd.n337 960
R2822 dvdd.n402 dvdd.n337 960
R2823 dvdd.n402 dvdd.n292 960
R2824 dvdd.n569 dvdd.n292 960
R2825 dvdd.n569 dvdd.n293 960
R2826 dvdd.n561 dvdd.n293 960
R2827 dvdd.n561 dvdd.n302 960
R2828 dvdd.n557 dvdd.n302 960
R2829 dvdd.n557 dvdd.n305 960
R2830 dvdd.n549 dvdd.n305 960
R2831 dvdd.n386 dvdd.n342 960
R2832 dvdd.n396 dvdd.n342 960
R2833 dvdd.n396 dvdd.n343 960
R2834 dvdd.n343 dvdd.n336 960
R2835 dvdd.n336 dvdd.n295 960
R2836 dvdd.n567 dvdd.n295 960
R2837 dvdd.n567 dvdd.n296 960
R2838 dvdd.n563 dvdd.n296 960
R2839 dvdd.n563 dvdd.n300 960
R2840 dvdd.n555 dvdd.n300 960
R2841 dvdd.n555 dvdd.n307 960
R2842 dvdd.n551 dvdd.n307 960
R2843 dvdd.n551 dvdd.n310 960
R2844 dvdd.n417 dvdd.n310 960
R2845 dvdd.n354 dvdd.n347 960
R2846 dvdd.n357 dvdd.n347 960
R2847 dvdd.n357 dvdd.n341 960
R2848 dvdd.n341 dvdd.n331 960
R2849 dvdd.n404 dvdd.n331 960
R2850 dvdd.n404 dvdd.n332 960
R2851 dvdd.n332 dvdd.n294 960
R2852 dvdd.n323 dvdd.n294 960
R2853 dvdd.n323 dvdd.n301 960
R2854 dvdd.n318 dvdd.n301 960
R2855 dvdd.n318 dvdd.n306 960
R2856 dvdd.n313 dvdd.n306 960
R2857 dvdd.n313 dvdd.n311 960
R2858 dvdd.n418 dvdd.n311 960
R2859 dvdd.n418 dvdd.n415 960
R2860 dvdd.n283 dvdd 925.605
R2861 dvdd.n354 dvdd.n346 878.823
R2862 dvdd.n358 dvdd.n357 878.823
R2863 dvdd.n358 dvdd.n342 878.823
R2864 dvdd.n391 dvdd.n331 878.823
R2865 dvdd.n391 dvdd.n343 878.823
R2866 dvdd.n333 dvdd.n332 878.823
R2867 dvdd.n333 dvdd.n295 878.823
R2868 dvdd.n324 dvdd.n323 878.823
R2869 dvdd.n324 dvdd.n296 878.823
R2870 dvdd.n321 dvdd.n318 878.823
R2871 dvdd.n321 dvdd.n300 878.823
R2872 dvdd.n418 dvdd.n312 878.823
R2873 dvdd.n316 dvdd.n305 878.823
R2874 dvdd.n316 dvdd.n313 878.823
R2875 dvdd.n319 dvdd.n302 878.823
R2876 dvdd.n319 dvdd.n318 878.823
R2877 dvdd.n326 dvdd.n293 878.823
R2878 dvdd.n326 dvdd.n323 878.823
R2879 dvdd.n334 dvdd.n292 878.823
R2880 dvdd.n334 dvdd.n332 878.823
R2881 dvdd.n389 dvdd.n337 878.823
R2882 dvdd.n389 dvdd.n331 878.823
R2883 dvdd.n360 dvdd.n340 878.823
R2884 dvdd.n360 dvdd.n357 878.823
R2885 dvdd.n353 dvdd.n348 878.823
R2886 dvdd.n354 dvdd.n353 878.823
R2887 dvdd.n314 dvdd.n313 878.823
R2888 dvdd.n314 dvdd.n307 878.823
R2889 dvdd.n420 dvdd.n418 878.823
R2890 dvdd.n420 dvdd.n310 878.823
R2891 dvdd.n377 dvdd.n355 878.823
R2892 dvdd.n368 dvdd.n351 878.823
R2893 dvdd.n170 dvdd.t2 869.832
R2894 dvdd.n229 dvdd.t109 856.909
R2895 dvdd.n260 dvdd.t1 848.84
R2896 dvdd.n380 dvdd.n348 818.823
R2897 dvdd.n370 dvdd.n355 818.823
R2898 dvdd.n151 dvdd.n146 772.942
R2899 dvdd.n151 dvdd.n148 772.942
R2900 dvdd.n594 dvdd.n583 741.178
R2901 dvdd.n612 dvdd.n583 741.178
R2902 dvdd.n612 dvdd.n584 741.178
R2903 dvdd.n596 dvdd.n590 741.178
R2904 dvdd.n590 dvdd.n585 741.178
R2905 dvdd.n586 dvdd.n585 741.178
R2906 dvdd.n453 dvdd.n446 741.178
R2907 dvdd.n451 dvdd.n442 741.178
R2908 dvdd.n153 dvdd.n146 741.178
R2909 dvdd.n161 dvdd.n146 741.178
R2910 dvdd.n155 dvdd.n148 741.178
R2911 dvdd.n159 dvdd.n148 741.178
R2912 dvdd.n201 dvdd.t330 685.053
R2913 dvdd.n222 dvdd.n186 682.808
R2914 dvdd.n239 dvdd.t328 680.702
R2915 dvdd.n238 dvdd.t326 674.558
R2916 dvdd.n236 dvdd.t218 667.346
R2917 dvdd.n266 dvdd.t210 661.764
R2918 dvdd.n265 dvdd.t208 661.663
R2919 dvdd.n188 dvdd.n187 611.958
R2920 dvdd.n505 dvdd.n493 610.588
R2921 dvdd.n505 dvdd.n504 610.588
R2922 dvdd.n498 dvdd.n494 610.588
R2923 dvdd.n508 dvdd.n498 610.588
R2924 dvdd.n208 dvdd.n207 610.407
R2925 dvdd.n193 dvdd.n192 607.497
R2926 dvdd.n181 dvdd.n180 606.721
R2927 dvdd.n101 dvdd.n97 604.213
R2928 dvdd.n116 dvdd.n110 604.213
R2929 dvdd.n231 dvdd.n183 601.292
R2930 dvdd.n247 dvdd.n176 597.51
R2931 dvdd.n602 dvdd.n584 557.648
R2932 dvdd.n605 dvdd.n586 557.648
R2933 dvdd.n530 dvdd.n446 557.648
R2934 dvdd.n530 dvdd.n447 557.648
R2935 dvdd.n526 dvdd.n447 557.648
R2936 dvdd.n526 dvdd.n461 557.648
R2937 dvdd.n490 dvdd.n461 557.648
R2938 dvdd.n531 dvdd.n442 557.648
R2939 dvdd.n531 dvdd.n443 557.648
R2940 dvdd.n462 dvdd.n443 557.648
R2941 dvdd.n463 dvdd.n462 557.648
R2942 dvdd.n520 dvdd.n463 557.648
R2943 dvdd.n101 dvdd.n96 556.98
R2944 dvdd.n110 dvdd.n108 556.819
R2945 dvdd dvdd.t65 516.562
R2946 dvdd.n370 dvdd.n368 465.882
R2947 dvdd dvdd.t211 415.625
R2948 dvdd.n282 dvdd 384.986
R2949 dvdd.n513 dvdd.n495 371.2
R2950 dvdd.n355 dvdd.n354 352.942
R2951 dvdd.n139 dvdd.t72 346.464
R2952 dvdd.n138 dvdd.t20 346.421
R2953 dvdd.n0 dvdd.t107 346.406
R2954 dvdd.n1 dvdd.t104 346.385
R2955 dvdd.n81 dvdd.t294 346.253
R2956 dvdd.n80 dvdd.t139 346.253
R2957 dvdd.n81 dvdd.t266 345.885
R2958 dvdd.n80 dvdd.t297 345.885
R2959 dvdd.n1 dvdd.t105 345.849
R2960 dvdd.n138 dvdd.t179 345.844
R2961 dvdd.n139 dvdd.t18 345.841
R2962 dvdd.n0 dvdd.t346 345.841
R2963 dvdd.n215 dvdd.t286 342.274
R2964 dvdd.n140 dvdd.t178 340.822
R2965 dvdd.n438 dvdd.t4 340.692
R2966 dvdd.n465 dvdd.t182 340.685
R2967 dvdd.n467 dvdd.t50 340.68
R2968 dvdd.n140 dvdd.t177 340.219
R2969 dvdd.n467 dvdd.t313 340.217
R2970 dvdd.n465 dvdd.t181 340.212
R2971 dvdd.n438 dvdd.t221 340.209
R2972 dvdd.n262 dvdd.n261 333.271
R2973 dvdd.t207 dvdd.n269 332.31
R2974 dvdd.t209 dvdd.n270 332.31
R2975 dvdd.n196 dvdd.n195 325.743
R2976 dvdd.n174 dvdd.n173 325.255
R2977 dvdd.n169 dvdd.n168 322.68
R2978 dvdd.n246 dvdd.n177 320.902
R2979 dvdd.n254 dvdd.n172 320.902
R2980 dvdd.n203 dvdd.n202 319.026
R2981 dvdd.n423 dvdd.t154 318.216
R2982 dvdd.n285 dvdd.t141 314.976
R2983 dvdd.n260 dvdd.t350 308.478
R2984 dvdd.t59 dvdd.n150 303.264
R2985 dvdd.t305 dvdd.n147 303.264
R2986 dvdd.n437 dvdd.n435 299.887
R2987 dvdd.n165 dvdd.n142 299.887
R2988 dvdd.n79 dvdd.n77 299.817
R2989 dvdd.n73 dvdd.n71 299.817
R2990 dvdd.n67 dvdd.n65 299.817
R2991 dvdd.n61 dvdd.n59 299.817
R2992 dvdd.n55 dvdd.n53 299.817
R2993 dvdd.n49 dvdd.n47 299.817
R2994 dvdd.n43 dvdd.n41 299.817
R2995 dvdd.n37 dvdd.n35 299.817
R2996 dvdd.n31 dvdd.n29 299.817
R2997 dvdd.n25 dvdd.n23 299.817
R2998 dvdd.n19 dvdd.n17 299.817
R2999 dvdd.n13 dvdd.n11 299.817
R3000 dvdd.n7 dvdd.n5 299.817
R3001 dvdd.n4 dvdd.n2 299.817
R3002 dvdd.n10 dvdd.n8 299.817
R3003 dvdd.n16 dvdd.n14 299.817
R3004 dvdd.n22 dvdd.n20 299.817
R3005 dvdd.n28 dvdd.n26 299.817
R3006 dvdd.n34 dvdd.n32 299.817
R3007 dvdd.n40 dvdd.n38 299.817
R3008 dvdd.n46 dvdd.n44 299.817
R3009 dvdd.n52 dvdd.n50 299.817
R3010 dvdd.n58 dvdd.n56 299.817
R3011 dvdd.n64 dvdd.n62 299.817
R3012 dvdd.n70 dvdd.n68 299.817
R3013 dvdd.n76 dvdd.n74 299.817
R3014 dvdd.n166 dvdd.n141 299.815
R3015 dvdd.n79 dvdd.n78 299.449
R3016 dvdd.n73 dvdd.n72 299.449
R3017 dvdd.n67 dvdd.n66 299.449
R3018 dvdd.n61 dvdd.n60 299.449
R3019 dvdd.n55 dvdd.n54 299.449
R3020 dvdd.n49 dvdd.n48 299.449
R3021 dvdd.n43 dvdd.n42 299.449
R3022 dvdd.n37 dvdd.n36 299.449
R3023 dvdd.n31 dvdd.n30 299.449
R3024 dvdd.n25 dvdd.n24 299.449
R3025 dvdd.n19 dvdd.n18 299.449
R3026 dvdd.n13 dvdd.n12 299.449
R3027 dvdd.n7 dvdd.n6 299.449
R3028 dvdd.n4 dvdd.n3 299.449
R3029 dvdd.n10 dvdd.n9 299.449
R3030 dvdd.n16 dvdd.n15 299.449
R3031 dvdd.n22 dvdd.n21 299.449
R3032 dvdd.n28 dvdd.n27 299.449
R3033 dvdd.n34 dvdd.n33 299.449
R3034 dvdd.n40 dvdd.n39 299.449
R3035 dvdd.n46 dvdd.n45 299.449
R3036 dvdd.n52 dvdd.n51 299.449
R3037 dvdd.n58 dvdd.n57 299.449
R3038 dvdd.n64 dvdd.n63 299.449
R3039 dvdd.n70 dvdd.n69 299.449
R3040 dvdd.n76 dvdd.n75 299.449
R3041 dvdd.n437 dvdd.n436 299.414
R3042 dvdd.n515 dvdd.n514 289.281
R3043 dvdd.t323 dvdd.n476 281.277
R3044 dvdd.n478 dvdd.t321 281.277
R3045 dvdd.t61 dvdd.n152 266.264
R3046 dvdd.n152 dvdd.t308 266.264
R3047 dvdd.n178 dvdd.t125 259.171
R3048 dvdd.n216 dvdd.t339 259.103
R3049 dvdd.n474 dvdd.n471 258.767
R3050 dvdd.t265 dvdd.n99 252.591
R3051 dvdd.t303 dvdd.n100 252.591
R3052 dvdd.t138 dvdd.n114 252.591
R3053 dvdd.n115 dvdd.t200 252.591
R3054 dvdd.t262 dvdd.n421 251.499
R3055 dvdd.n167 dvdd.t243 250.96
R3056 dvdd.n255 dvdd.t348 248.715
R3057 dvdd.n503 dvdd.n497 241.386
R3058 dvdd.n597 dvdd.n588 232.282
R3059 dvdd.n454 dvdd.n448 232.282
R3060 dvdd.n104 dvdd.n98 231.615
R3061 dvdd.n113 dvdd.n109 231.615
R3062 dvdd.n468 dvdd.t175 231.103
R3063 dvdd.n425 dvdd.t300 230.934
R3064 dvdd.n542 dvdd.t272 230.873
R3065 dvdd.n541 dvdd.t157 230.847
R3066 dvdd.n540 dvdd.t86 230.845
R3067 dvdd.n538 dvdd.t267 230.82
R3068 dvdd.n539 dvdd.t279 230.819
R3069 dvdd.n536 dvdd.t152 230.817
R3070 dvdd.n573 dvdd.t117 230.815
R3071 dvdd.n574 dvdd.t302 230.808
R3072 dvdd.n537 dvdd.t56 230.803
R3073 dvdd.n289 dvdd.t44 230.8
R3074 dvdd.n544 dvdd.t155 230.751
R3075 dvdd.n433 dvdd.t34 230.712
R3076 dvdd.n434 dvdd.t263 230.709
R3077 dvdd.n432 dvdd.t254 230.692
R3078 dvdd.n427 dvdd.t166 230.691
R3079 dvdd.n425 dvdd.t165 230.69
R3080 dvdd.n430 dvdd.t185 230.69
R3081 dvdd.n431 dvdd.t41 230.689
R3082 dvdd.n429 dvdd.t145 230.681
R3083 dvdd.n426 dvdd.t143 230.681
R3084 dvdd.n428 dvdd.t298 230.68
R3085 dvdd.n577 dvdd.t288 230.679
R3086 dvdd.n576 dvdd.t290 230.632
R3087 dvdd.n484 dvdd.t336 230.613
R3088 dvdd.n468 dvdd.t316 230.47
R3089 dvdd.n485 dvdd.t337 230.468
R3090 dvdd.t331 dvdd.t252 226.124
R3091 dvdd.n475 dvdd.t324 222.696
R3092 dvdd.n470 dvdd.t322 222.696
R3093 dvdd.n501 dvdd.n495 218.894
R3094 dvdd.n606 dvdd.n600 212.713
R3095 dvdd.n492 dvdd.n491 212.707
R3096 dvdd.n283 dvdd.t108 211.881
R3097 dvdd.n281 dvdd.n169 211.838
R3098 dvdd.n280 dvdd.n279 208.21
R3099 dvdd.n575 dvdd.n288 202.185
R3100 dvdd.n509 dvdd.n497 200.804
R3101 dvdd.n387 dvdd.n345 196.142
R3102 dvdd.n546 dvdd.n424 196.142
R3103 dvdd.n424 dvdd.n416 196.142
R3104 dvdd.n475 dvdd.n474 192.24
R3105 dvdd.n375 dvdd.n374 181.083
R3106 dvdd.n376 dvdd.n375 181.083
R3107 dvdd.t103 dvdd.n589 179.821
R3108 dvdd.t273 dvdd.n449 179.821
R3109 dvdd.n502 dvdd.n496 175.812
R3110 dvdd.n510 dvdd.n496 175.435
R3111 dvdd.n517 dvdd.t174 172.275
R3112 dvdd.n507 dvdd.t174 172.275
R3113 dvdd.n507 dvdd.t335 172.275
R3114 dvdd.n500 dvdd.n499 169.032
R3115 dvdd.n593 dvdd.n588 165.964
R3116 dvdd.n450 dvdd.n448 165.409
R3117 dvdd.n601 dvdd.n600 163.114
R3118 dvdd.n158 dvdd.n145 161.506
R3119 dvdd.n156 dvdd.n149 161.506
R3120 dvdd.t106 dvdd.n592 161.321
R3121 dvdd.n592 dvdd.t19 161.321
R3122 dvdd.t17 dvdd.n610 161.321
R3123 dvdd.t275 dvdd.n444 161.321
R3124 dvdd.n610 dvdd.t176 157.339
R3125 dvdd.t3 dvdd.n444 157.339
R3126 dvdd.t3 dvdd.n445 157.339
R3127 dvdd.t180 dvdd.n445 157.339
R3128 dvdd.t180 dvdd.n525 157.339
R3129 dvdd.n525 dvdd.t49 157.339
R3130 dvdd.n518 dvdd.t49 157.339
R3131 dvdd.n352 dvdd.t14 156.709
R3132 dvdd.n359 dvdd.t12 156.709
R3133 dvdd.n359 dvdd.t13 156.709
R3134 dvdd.n390 dvdd.t11 156.709
R3135 dvdd.n390 dvdd.t299 156.709
R3136 dvdd.t116 dvdd.n335 156.709
R3137 dvdd.n335 dvdd.t43 156.709
R3138 dvdd.n325 dvdd.t151 156.709
R3139 dvdd.n325 dvdd.t55 156.709
R3140 dvdd.n320 dvdd.t144 156.709
R3141 dvdd.n320 dvdd.t184 156.709
R3142 dvdd.n315 dvdd.t40 156.709
R3143 dvdd.n315 dvdd.t156 156.709
R3144 dvdd.n421 dvdd.t33 156.709
R3145 dvdd dvdd.t124 156.438
R3146 dvdd.n604 dvdd.n603 154.983
R3147 dvdd.n271 dvdd.n268 153.976
R3148 dvdd.n271 dvdd.n267 153.976
R3149 dvdd.n608 dvdd.n582 153.225
R3150 dvdd.n608 dvdd.n607 153.225
R3151 dvdd.n587 dvdd.n581 153.225
R3152 dvdd.n598 dvdd.n587 153.225
R3153 dvdd.n523 dvdd.n460 153.225
R3154 dvdd.n528 dvdd.n459 153.225
R3155 dvdd.n457 dvdd.n456 153.225
R3156 dvdd.n512 dvdd.n492 152.847
R3157 dvdd.n523 dvdd.n522 152.847
R3158 dvdd.n459 dvdd.n441 152.847
R3159 dvdd.n456 dvdd.n440 152.847
R3160 dvdd.n180 dvdd.t161 150.827
R3161 dvdd.n373 dvdd.n372 143.852
R3162 dvdd.t130 dvdd.t132 142.216
R3163 dvdd.t327 dvdd 140.793
R3164 dvdd.n284 dvdd 139.531
R3165 dvdd.t242 dvdd.t331 139.371
R3166 dvdd.t0 dvdd 136.528
R3167 dvdd.t219 dvdd.t203 132.024
R3168 dvdd.t292 dvdd.t265 131.412
R3169 dvdd.t98 dvdd.t292 131.412
R3170 dvdd.t38 dvdd.t98 131.412
R3171 dvdd.t31 dvdd.t38 131.412
R3172 dvdd.t162 dvdd.t31 131.412
R3173 dvdd.t5 dvdd.t162 131.412
R3174 dvdd.t45 dvdd.t5 131.412
R3175 dvdd.t73 dvdd.t45 131.412
R3176 dvdd.t268 dvdd.t73 131.412
R3177 dvdd.t7 dvdd.t268 131.412
R3178 dvdd.t100 dvdd.t7 131.412
R3179 dvdd.t29 dvdd.t100 131.412
R3180 dvdd.t96 dvdd.t29 131.412
R3181 dvdd.t96 dvdd.t47 131.412
R3182 dvdd.t47 dvdd.t57 131.412
R3183 dvdd.t57 dvdd.t311 131.412
R3184 dvdd.t311 dvdd.t205 131.412
R3185 dvdd.t205 dvdd.t77 131.412
R3186 dvdd.t77 dvdd.t27 131.412
R3187 dvdd.t27 dvdd.t192 131.412
R3188 dvdd.t192 dvdd.t23 131.412
R3189 dvdd.t23 dvdd.t21 131.412
R3190 dvdd.t21 dvdd.t25 131.412
R3191 dvdd.t25 dvdd.t186 131.412
R3192 dvdd.t186 dvdd.t188 131.412
R3193 dvdd.t188 dvdd.t303 131.412
R3194 dvdd.t70 dvdd.t138 131.412
R3195 dvdd.t255 dvdd.t70 131.412
R3196 dvdd.t53 dvdd.t255 131.412
R3197 dvdd.t259 dvdd.t53 131.412
R3198 dvdd.t51 dvdd.t259 131.412
R3199 dvdd.t270 dvdd.t51 131.412
R3200 dvdd.t112 dvdd.t270 131.412
R3201 dvdd.t146 dvdd.t112 131.412
R3202 dvdd.t257 dvdd.t146 131.412
R3203 dvdd.t79 dvdd.t257 131.412
R3204 dvdd.t82 dvdd.t79 131.412
R3205 dvdd.t195 dvdd.t82 131.412
R3206 dvdd.t148 dvdd.t195 131.412
R3207 dvdd.t84 dvdd.t148 131.412
R3208 dvdd.t295 dvdd.t84 131.412
R3209 dvdd.t227 dvdd.t295 131.412
R3210 dvdd.t63 dvdd.t227 131.412
R3211 dvdd.t94 dvdd.t63 131.412
R3212 dvdd.t224 dvdd.t94 131.412
R3213 dvdd.t92 dvdd.t224 131.412
R3214 dvdd.t229 dvdd.t92 131.412
R3215 dvdd.t231 dvdd.t229 131.412
R3216 dvdd.t90 dvdd.t231 131.412
R3217 dvdd.t280 dvdd.t90 131.412
R3218 dvdd.t283 dvdd.t280 131.412
R3219 dvdd.t200 dvdd.t283 131.412
R3220 dvdd.n374 dvdd.n367 131.338
R3221 dvdd.t36 dvdd.t160 130.175
R3222 dvdd.t246 dvdd.t244 127.995
R3223 dvdd.t244 dvdd.t248 127.995
R3224 dvdd.t122 dvdd 125.15
R3225 dvdd.t212 dvdd.t36 124.636
R3226 dvdd.n282 dvdd.t171 123.156
R3227 dvdd.t217 dvdd.t325 122.305
R3228 dvdd.t164 dvdd.t134 122.305
R3229 dvdd dvdd.t169 121.98
R3230 dvdd.n548 dvdd.n547 121.156
R3231 dvdd.t75 dvdd.t126 118.04
R3232 dvdd.n381 dvdd.n350 117.93
R3233 dvdd.n422 dvdd.t262 117.633
R3234 dvdd.t154 dvdd.n422 117.633
R3235 dvdd.n192 dvdd.t10 112.572
R3236 dvdd.t120 dvdd.t67 112.35
R3237 dvdd.t110 dvdd.t223 112.35
R3238 dvdd.n202 dvdd.t251 110.227
R3239 dvdd.n186 dvdd.t220 110.227
R3240 dvdd.n186 dvdd.t16 110.227
R3241 dvdd.n518 dvdd.n517 105.556
R3242 dvdd.n388 dvdd.n387 102.4
R3243 dvdd.n395 dvdd.n388 102.4
R3244 dvdd.n395 dvdd.n394 102.4
R3245 dvdd.n394 dvdd.n393 102.4
R3246 dvdd.n393 dvdd.n297 102.4
R3247 dvdd.n566 dvdd.n297 102.4
R3248 dvdd.n566 dvdd.n565 102.4
R3249 dvdd.n565 dvdd.n564 102.4
R3250 dvdd.n564 dvdd.n299 102.4
R3251 dvdd.n554 dvdd.n299 102.4
R3252 dvdd.n554 dvdd.n553 102.4
R3253 dvdd.n553 dvdd.n552 102.4
R3254 dvdd.n552 dvdd.n309 102.4
R3255 dvdd.n416 dvdd.n309 102.4
R3256 dvdd.n365 dvdd.n364 102.4
R3257 dvdd.n364 dvdd.n363 102.4
R3258 dvdd.n363 dvdd.n362 102.4
R3259 dvdd.n362 dvdd.n330 102.4
R3260 dvdd.n405 dvdd.n330 102.4
R3261 dvdd.n406 dvdd.n405 102.4
R3262 dvdd.n407 dvdd.n406 102.4
R3263 dvdd.n408 dvdd.n407 102.4
R3264 dvdd.n409 dvdd.n408 102.4
R3265 dvdd.n410 dvdd.n409 102.4
R3266 dvdd.n411 dvdd.n410 102.4
R3267 dvdd.n412 dvdd.n411 102.4
R3268 dvdd.n413 dvdd.n412 102.4
R3269 dvdd.n414 dvdd.n413 102.4
R3270 dvdd.n546 dvdd.n414 102.4
R3271 dvdd.t329 dvdd.t250 102.395
R3272 dvdd.t9 dvdd.t215 102.395
R3273 dvdd.n207 dvdd.t216 100.846
R3274 dvdd.n207 dvdd.t68 98.5005
R3275 dvdd.t223 dvdd.n284 98.1292
R3276 dvdd.n547 dvdd.n546 97.7422
R3277 dvdd.n477 dvdd.t323 94.5219
R3278 dvdd.t321 dvdd.n477 94.5219
R3279 dvdd.n365 dvdd.n345 93.7417
R3280 dvdd.n363 dvdd.n344 93.7417
R3281 dvdd.n388 dvdd.n344 93.7417
R3282 dvdd.n361 dvdd.n339 93.7417
R3283 dvdd.n363 dvdd.n361 93.7417
R3284 dvdd.n392 dvdd.n330 93.7417
R3285 dvdd.n394 dvdd.n392 93.7417
R3286 dvdd.n400 dvdd.n338 93.7417
R3287 dvdd.n338 dvdd.n330 93.7417
R3288 dvdd.n406 dvdd.n328 93.7417
R3289 dvdd.n328 dvdd.n297 93.7417
R3290 dvdd.n329 dvdd.n290 93.7417
R3291 dvdd.n406 dvdd.n329 93.7417
R3292 dvdd.n408 dvdd.n298 93.7417
R3293 dvdd.n565 dvdd.n298 93.7417
R3294 dvdd.n327 dvdd.n291 93.7417
R3295 dvdd.n408 dvdd.n327 93.7417
R3296 dvdd.n410 dvdd.n322 93.7417
R3297 dvdd.n322 dvdd.n299 93.7417
R3298 dvdd.n559 dvdd.n303 93.7417
R3299 dvdd.n410 dvdd.n303 93.7417
R3300 dvdd.n317 dvdd.n304 93.7417
R3301 dvdd.n412 dvdd.n317 93.7417
R3302 dvdd.n382 dvdd.n349 93.7417
R3303 dvdd.n365 dvdd.n349 93.7417
R3304 dvdd.n412 dvdd.n308 93.7417
R3305 dvdd.n553 dvdd.n308 93.7417
R3306 dvdd.n419 dvdd.n414 93.7417
R3307 dvdd.n419 dvdd.n309 93.7417
R3308 dvdd.n376 dvdd.n366 93.7417
R3309 dvdd.n367 dvdd.n350 92.8212
R3310 dvdd.n606 dvdd.n605 92.5005
R3311 dvdd.n602 dvdd.n601 92.5005
R3312 dvdd.n602 dvdd.t176 92.5005
R3313 dvdd.n530 dvdd.n529 92.5005
R3314 dvdd.t3 dvdd.n530 92.5005
R3315 dvdd.n527 dvdd.n526 92.5005
R3316 dvdd.n526 dvdd.t180 92.5005
R3317 dvdd.n491 dvdd.n490 92.5005
R3318 dvdd.n490 dvdd.t49 92.5005
R3319 dvdd.n521 dvdd.n520 92.5005
R3320 dvdd.n520 dvdd.t49 92.5005
R3321 dvdd.n464 dvdd.n462 92.5005
R3322 dvdd.t180 dvdd.n462 92.5005
R3323 dvdd.n532 dvdd.n531 92.5005
R3324 dvdd.n531 dvdd.t3 92.5005
R3325 dvdd.n162 dvdd.n145 91.8757
R3326 dvdd.n149 dvdd.n143 91.8757
R3327 dvdd.n275 dvdd.n268 91.6804
R3328 dvdd.n276 dvdd.n267 91.4705
R3329 dvdd.n187 dvdd.t170 91.4648
R3330 dvdd.t211 dvdd.t338 89.063
R3331 dvdd.n369 dvdd.n366 87.3417
R3332 dvdd.n273 dvdd.t207 84.7589
R3333 dvdd.n273 dvdd.t209 84.7589
R3334 dvdd.t240 dvdd.t130 83.9077
R3335 dvdd.t214 dvdd.t111 83.2331
R3336 dvdd.n157 dvdd.n144 82.4476
R3337 dvdd.n605 dvdd.n604 81.5301
R3338 dvdd.n378 dvdd.n352 81.1971
R3339 dvdd.n180 dvdd.t172 80.821
R3340 dvdd.n163 dvdd.n144 80.1887
R3341 dvdd.n598 dvdd.n597 79.0593
R3342 dvdd.n599 dvdd.n598 79.0593
R3343 dvdd.n607 dvdd.n599 79.0593
R3344 dvdd.n457 dvdd.n454 79.0593
R3345 dvdd.n157 dvdd.n156 79.0593
R3346 dvdd.n158 dvdd.n157 79.0593
R3347 dvdd.n154 dvdd.t59 78.8932
R3348 dvdd.n154 dvdd.t61 78.8932
R3349 dvdd.n160 dvdd.t308 78.8932
R3350 dvdd.n160 dvdd.t305 78.8932
R3351 dvdd.t347 dvdd.t122 78.2191
R3352 dvdd.n281 dvdd.t246 76.7969
R3353 dvdd.t132 dvdd.t35 72.5304
R3354 dvdd.n192 dvdd.t121 70.3576
R3355 dvdd.n187 dvdd.t204 70.3576
R3356 dvdd dvdd.n280 68.264
R3357 dvdd.n280 dvdd 68.264
R3358 dvdd.t15 dvdd.t66 66.0126
R3359 dvdd.n502 dvdd.n501 65.1299
R3360 dvdd.n503 dvdd.n502 65.1299
R3361 dvdd.n385 dvdd.t14 64.1458
R3362 dvdd.n385 dvdd.t12 64.1458
R3363 dvdd.n397 dvdd.t13 64.1458
R3364 dvdd.n397 dvdd.t11 64.1458
R3365 dvdd.n403 dvdd.t299 64.1458
R3366 dvdd.n403 dvdd.t116 64.1458
R3367 dvdd.n568 dvdd.t43 64.1458
R3368 dvdd.n568 dvdd.t151 64.1458
R3369 dvdd.n562 dvdd.t55 64.1458
R3370 dvdd.n562 dvdd.t144 64.1458
R3371 dvdd.n556 dvdd.t184 64.1458
R3372 dvdd.n556 dvdd.t40 64.1458
R3373 dvdd.n550 dvdd.t156 64.1458
R3374 dvdd.n550 dvdd.t33 64.1458
R3375 dvdd.t136 dvdd.t347 63.9975
R3376 dvdd.n509 dvdd.n508 61.6672
R3377 dvdd.n511 dvdd.n494 61.6672
R3378 dvdd.n501 dvdd.n493 61.6672
R3379 dvdd.n493 dvdd.t174 61.6672
R3380 dvdd.n504 dvdd.n503 61.6672
R3381 dvdd.n514 dvdd.n511 60.1048
R3382 dvdd.n607 dvdd.n606 59.4829
R3383 dvdd.n529 dvdd.n457 59.4829
R3384 dvdd.n529 dvdd.n528 59.4829
R3385 dvdd.n528 dvdd.n527 59.4829
R3386 dvdd.n527 dvdd.n460 59.4829
R3387 dvdd.n491 dvdd.n460 59.4829
R3388 dvdd.n372 dvdd.t317 59.274
R3389 dvdd.t289 dvdd.n378 59.274
R3390 dvdd.n471 dvdd.n470 55.9243
R3391 dvdd.n504 dvdd.n500 55.5369
R3392 dvdd.t35 dvdd.t136 55.4646
R3393 dvdd.t215 dvdd.t120 51.1981
R3394 dvdd.t128 dvdd.n281 51.1981
R3395 dvdd.t222 dvdd.n283 50.2271
R3396 dvdd.t252 dvdd.t329 49.7759
R3397 dvdd.n369 dvdd.n367 49.684
R3398 dvdd.t317 dvdd.n371 47.9065
R3399 dvdd.n379 dvdd.t289 47.9065
R3400 dvdd.n595 dvdd.t103 47.7992
R3401 dvdd.n595 dvdd.t106 47.7992
R3402 dvdd.n611 dvdd.t19 47.7992
R3403 dvdd.n611 dvdd.t17 47.7992
R3404 dvdd.n452 dvdd.t273 47.7992
R3405 dvdd.n452 dvdd.t275 47.7992
R3406 dvdd.n195 dvdd.t332 46.9053
R3407 dvdd.n435 dvdd.t274 46.4362
R3408 dvdd.n435 dvdd.t277 46.4362
R3409 dvdd.n436 dvdd.t278 46.4362
R3410 dvdd.n436 dvdd.t276 46.4362
R3411 dvdd.n141 dvdd.t309 46.4362
R3412 dvdd.n141 dvdd.t306 46.4362
R3413 dvdd.n142 dvdd.t60 46.4362
R3414 dvdd.n142 dvdd.t62 46.4362
R3415 dvdd.n77 dvdd.t293 46.4362
R3416 dvdd.n77 dvdd.t159 46.4362
R3417 dvdd.n78 dvdd.t344 46.4362
R3418 dvdd.n78 dvdd.t99 46.4362
R3419 dvdd.n71 dvdd.t39 46.4362
R3420 dvdd.n71 dvdd.t264 46.4362
R3421 dvdd.n72 dvdd.t102 46.4362
R3422 dvdd.n72 dvdd.t32 46.4362
R3423 dvdd.n65 dvdd.t163 46.4362
R3424 dvdd.n65 dvdd.t88 46.4362
R3425 dvdd.n66 dvdd.t183 46.4362
R3426 dvdd.n66 dvdd.t6 46.4362
R3427 dvdd.n59 dvdd.t46 46.4362
R3428 dvdd.n59 dvdd.t74 46.4362
R3429 dvdd.n60 dvdd.t87 46.4362
R3430 dvdd.n60 dvdd.t167 46.4362
R3431 dvdd.n53 dvdd.t343 46.4362
R3432 dvdd.n53 dvdd.t89 46.4362
R3433 dvdd.n54 dvdd.t269 46.4362
R3434 dvdd.n54 dvdd.t8 46.4362
R3435 dvdd.n47 dvdd.t101 46.4362
R3436 dvdd.n47 dvdd.t30 46.4362
R3437 dvdd.n48 dvdd.t114 46.4362
R3438 dvdd.n48 dvdd.t168 46.4362
R3439 dvdd.n41 dvdd.t97 46.4362
R3440 dvdd.n41 dvdd.t48 46.4362
R3441 dvdd.n42 dvdd.t291 46.4362
R3442 dvdd.n42 dvdd.t158 46.4362
R3443 dvdd.n35 dvdd.t58 46.4362
R3444 dvdd.n35 dvdd.t341 46.4362
R3445 dvdd.n36 dvdd.t115 46.4362
R3446 dvdd.n36 dvdd.t312 46.4362
R3447 dvdd.n29 dvdd.t206 46.4362
R3448 dvdd.n29 dvdd.t345 46.4362
R3449 dvdd.n30 dvdd.t340 46.4362
R3450 dvdd.n30 dvdd.t78 46.4362
R3451 dvdd.n23 dvdd.t315 46.4362
R3452 dvdd.n23 dvdd.t193 46.4362
R3453 dvdd.n24 dvdd.t28 46.4362
R3454 dvdd.n24 dvdd.t314 46.4362
R3455 dvdd.n17 dvdd.t24 46.4362
R3456 dvdd.n17 dvdd.t173 46.4362
R3457 dvdd.n18 dvdd.t194 46.4362
R3458 dvdd.n18 dvdd.t22 46.4362
R3459 dvdd.n11 dvdd.t26 46.4362
R3460 dvdd.n11 dvdd.t187 46.4362
R3461 dvdd.n12 dvdd.t310 46.4362
R3462 dvdd.n12 dvdd.t190 46.4362
R3463 dvdd.n5 dvdd.t191 46.4362
R3464 dvdd.n5 dvdd.t307 46.4362
R3465 dvdd.n6 dvdd.t189 46.4362
R3466 dvdd.n6 dvdd.t304 46.4362
R3467 dvdd.n3 dvdd.t284 46.4362
R3468 dvdd.n3 dvdd.t201 46.4362
R3469 dvdd.n2 dvdd.t285 46.4362
R3470 dvdd.n2 dvdd.t202 46.4362
R3471 dvdd.n9 dvdd.t236 46.4362
R3472 dvdd.n9 dvdd.t281 46.4362
R3473 dvdd.n8 dvdd.t91 46.4362
R3474 dvdd.n8 dvdd.t282 46.4362
R3475 dvdd.n15 dvdd.t230 46.4362
R3476 dvdd.n15 dvdd.t239 46.4362
R3477 dvdd.n14 dvdd.t237 46.4362
R3478 dvdd.n14 dvdd.t232 46.4362
R3479 dvdd.n21 dvdd.t233 46.4362
R3480 dvdd.n21 dvdd.t93 46.4362
R3481 dvdd.n20 dvdd.t225 46.4362
R3482 dvdd.n20 dvdd.t235 46.4362
R3483 dvdd.n27 dvdd.t226 46.4362
R3484 dvdd.n27 dvdd.t238 46.4362
R3485 dvdd.n26 dvdd.t64 46.4362
R3486 dvdd.n26 dvdd.t95 46.4362
R3487 dvdd.n33 dvdd.t333 46.4362
R3488 dvdd.n33 dvdd.t234 46.4362
R3489 dvdd.n32 dvdd.t296 46.4362
R3490 dvdd.n32 dvdd.t228 46.4362
R3491 dvdd.n39 dvdd.t149 46.4362
R3492 dvdd.n39 dvdd.t140 46.4362
R3493 dvdd.n38 dvdd.t334 46.4362
R3494 dvdd.n38 dvdd.t85 46.4362
R3495 dvdd.n45 dvdd.t83 46.4362
R3496 dvdd.n45 dvdd.t199 46.4362
R3497 dvdd.n44 dvdd.t150 46.4362
R3498 dvdd.n44 dvdd.t196 46.4362
R3499 dvdd.n51 dvdd.t258 46.4362
R3500 dvdd.n51 dvdd.t197 46.4362
R3501 dvdd.n50 dvdd.t301 46.4362
R3502 dvdd.n50 dvdd.t80 46.4362
R3503 dvdd.n57 dvdd.t113 46.4362
R3504 dvdd.n57 dvdd.t147 46.4362
R3505 dvdd.n56 dvdd.t342 46.4362
R3506 dvdd.n56 dvdd.t198 46.4362
R3507 dvdd.n63 dvdd.t52 46.4362
R3508 dvdd.n63 dvdd.t318 46.4362
R3509 dvdd.n62 dvdd.t81 46.4362
R3510 dvdd.n62 dvdd.t271 46.4362
R3511 dvdd.n69 dvdd.t69 46.4362
R3512 dvdd.n69 dvdd.t260 46.4362
R3513 dvdd.n68 dvdd.t54 46.4362
R3514 dvdd.n68 dvdd.t319 46.4362
R3515 dvdd.n75 dvdd.t153 46.4362
R3516 dvdd.n75 dvdd.t256 46.4362
R3517 dvdd.n74 dvdd.t71 46.4362
R3518 dvdd.n74 dvdd.t261 46.4362
R3519 dvdd.n599 dvdd.n585 46.2505
R3520 dvdd.n611 dvdd.n585 46.2505
R3521 dvdd.n597 dvdd.n596 46.2505
R3522 dvdd.n596 dvdd.n595 46.2505
R3523 dvdd.n594 dvdd.n593 46.2505
R3524 dvdd.n595 dvdd.n594 46.2505
R3525 dvdd.n613 dvdd.n612 46.2505
R3526 dvdd.n612 dvdd.n611 46.2505
R3527 dvdd.n454 dvdd.n453 46.2505
R3528 dvdd.n453 dvdd.n452 46.2505
R3529 dvdd.n451 dvdd.n450 46.2505
R3530 dvdd.n452 dvdd.n451 46.2505
R3531 dvdd.n270 dvdd.n268 46.2505
R3532 dvdd.n272 dvdd.n271 46.2505
R3533 dvdd.n273 dvdd.n272 46.2505
R3534 dvdd.n269 dvdd.n267 46.2505
R3535 dvdd.n275 dvdd.n274 46.2505
R3536 dvdd.n274 dvdd.n273 46.2505
R3537 dvdd.n159 dvdd.n158 46.2505
R3538 dvdd.n160 dvdd.n159 46.2505
R3539 dvdd.n156 dvdd.n155 46.2505
R3540 dvdd.n155 dvdd.n154 46.2505
R3541 dvdd.n153 dvdd.n143 46.2505
R3542 dvdd.n154 dvdd.n153 46.2505
R3543 dvdd.n162 dvdd.n161 46.2505
R3544 dvdd.n161 dvdd.n160 46.2505
R3545 dvdd.t203 dvdd.t15 45.9219
R3546 dvdd.t66 dvdd.t214 45.9219
R3547 dvdd.t111 dvdd.t222 45.9219
R3548 dvdd.t126 dvdd.t240 44.0873
R3549 dvdd.n515 dvdd.n495 38.4005
R3550 dvdd.n176 dvdd.t241 37.8175
R3551 dvdd.n366 dvdd.n365 37.6476
R3552 dvdd.n381 dvdd.n380 37.0005
R3553 dvdd.n380 dvdd.n379 37.0005
R3554 dvdd.n375 dvdd.n356 37.0005
R3555 dvdd.n371 dvdd.n356 37.0005
R3556 dvdd.n370 dvdd.n369 37.0005
R3557 dvdd.n371 dvdd.n370 37.0005
R3558 dvdd.n151 dvdd.n144 37.0005
R3559 dvdd.n152 dvdd.n151 37.0005
R3560 dvdd.n147 dvdd.n145 37.0005
R3561 dvdd.n150 dvdd.n149 37.0005
R3562 dvdd.n210 dvdd.n209 36.1417
R3563 dvdd.n210 dvdd.n190 36.1417
R3564 dvdd.n214 dvdd.n190 36.1417
R3565 dvdd.n218 dvdd.n217 36.1417
R3566 dvdd.n224 dvdd.n223 36.1417
R3567 dvdd.n224 dvdd.n184 36.1417
R3568 dvdd.n228 dvdd.n184 36.1417
R3569 dvdd.n245 dvdd.n244 36.1417
R3570 dvdd.n253 dvdd.n252 36.1417
R3571 dvdd.n176 dvdd.t76 36.0585
R3572 dvdd.n232 dvdd.n181 35.7652
R3573 dvdd.n223 dvdd.n222 35.3887
R3574 dvdd.n232 dvdd.n231 35.3887
R3575 dvdd.n202 dvdd.t253 35.1791
R3576 dvdd.n173 dvdd.t131 35.1791
R3577 dvdd.n172 dvdd.t137 35.1791
R3578 dvdd.n238 dvdd.n237 33.5064
R3579 dvdd.n475 dvdd.n469 33.4576
R3580 dvdd.n371 dvdd.t287 33.2911
R3581 dvdd.n379 dvdd.t320 33.2911
R3582 dvdd.n177 dvdd.t135 32.5407
R3583 dvdd.n195 dvdd.t142 32.1717
R3584 dvdd.n237 dvdd.n236 32.0005
R3585 dvdd.n218 dvdd.n188 31.2476
R3586 dvdd.n99 dvdd.n98 30.8338
R3587 dvdd.n100 dvdd.n97 30.8338
R3588 dvdd.n116 dvdd.n115 30.8338
R3589 dvdd.n114 dvdd.n113 30.8338
R3590 dvdd.n353 dvdd.n349 30.8338
R3591 dvdd.n353 dvdd.n352 30.8338
R3592 dvdd.n547 dvdd.n312 30.8338
R3593 dvdd.n421 dvdd.n312 30.8338
R3594 dvdd.n317 dvdd.n316 30.8338
R3595 dvdd.n316 dvdd.n315 30.8338
R3596 dvdd.n319 dvdd.n303 30.8338
R3597 dvdd.n320 dvdd.n319 30.8338
R3598 dvdd.n322 dvdd.n321 30.8338
R3599 dvdd.n321 dvdd.n320 30.8338
R3600 dvdd.n327 dvdd.n326 30.8338
R3601 dvdd.n326 dvdd.n325 30.8338
R3602 dvdd.n324 dvdd.n298 30.8338
R3603 dvdd.n325 dvdd.n324 30.8338
R3604 dvdd.n334 dvdd.n329 30.8338
R3605 dvdd.n335 dvdd.n334 30.8338
R3606 dvdd.n333 dvdd.n328 30.8338
R3607 dvdd.n335 dvdd.n333 30.8338
R3608 dvdd.n389 dvdd.n338 30.8338
R3609 dvdd.n390 dvdd.n389 30.8338
R3610 dvdd.n392 dvdd.n391 30.8338
R3611 dvdd.n391 dvdd.n390 30.8338
R3612 dvdd.n361 dvdd.n360 30.8338
R3613 dvdd.n360 dvdd.n359 30.8338
R3614 dvdd.n358 dvdd.n344 30.8338
R3615 dvdd.n359 dvdd.n358 30.8338
R3616 dvdd.n346 dvdd.n345 30.8338
R3617 dvdd.n352 dvdd.n346 30.8338
R3618 dvdd.n314 dvdd.n308 30.8338
R3619 dvdd.n315 dvdd.n314 30.8338
R3620 dvdd.n420 dvdd.n419 30.8338
R3621 dvdd.n421 dvdd.n420 30.8338
R3622 dvdd.n417 dvdd.n416 30.8338
R3623 dvdd.n422 dvdd.n417 30.8338
R3624 dvdd.n552 dvdd.n551 30.8338
R3625 dvdd.n551 dvdd.n550 30.8338
R3626 dvdd.n555 dvdd.n554 30.8338
R3627 dvdd.n556 dvdd.n555 30.8338
R3628 dvdd.n564 dvdd.n563 30.8338
R3629 dvdd.n563 dvdd.n562 30.8338
R3630 dvdd.n567 dvdd.n566 30.8338
R3631 dvdd.n568 dvdd.n567 30.8338
R3632 dvdd.n393 dvdd.n336 30.8338
R3633 dvdd.n403 dvdd.n336 30.8338
R3634 dvdd.n396 dvdd.n395 30.8338
R3635 dvdd.n397 dvdd.n396 30.8338
R3636 dvdd.n387 dvdd.n386 30.8338
R3637 dvdd.n386 dvdd.n385 30.8338
R3638 dvdd.n424 dvdd.n423 30.8338
R3639 dvdd.n351 dvdd.n350 30.8338
R3640 dvdd.n372 dvdd.n351 30.8338
R3641 dvdd.n384 dvdd.n383 30.8338
R3642 dvdd.n385 dvdd.n384 30.8338
R3643 dvdd.n399 dvdd.n398 30.8338
R3644 dvdd.n398 dvdd.n397 30.8338
R3645 dvdd.n402 dvdd.n401 30.8338
R3646 dvdd.n403 dvdd.n402 30.8338
R3647 dvdd.n570 dvdd.n569 30.8338
R3648 dvdd.n569 dvdd.n568 30.8338
R3649 dvdd.n561 dvdd.n560 30.8338
R3650 dvdd.n562 dvdd.n561 30.8338
R3651 dvdd.n558 dvdd.n557 30.8338
R3652 dvdd.n557 dvdd.n556 30.8338
R3653 dvdd.n549 dvdd.n548 30.8338
R3654 dvdd.n550 dvdd.n549 30.8338
R3655 dvdd.n374 dvdd.n373 30.8338
R3656 dvdd.n377 dvdd.n376 30.8338
R3657 dvdd.n378 dvdd.n377 30.8338
R3658 dvdd.n364 dvdd.n347 30.8338
R3659 dvdd.n385 dvdd.n347 30.8338
R3660 dvdd.n362 dvdd.n341 30.8338
R3661 dvdd.n397 dvdd.n341 30.8338
R3662 dvdd.n405 dvdd.n404 30.8338
R3663 dvdd.n404 dvdd.n403 30.8338
R3664 dvdd.n407 dvdd.n294 30.8338
R3665 dvdd.n568 dvdd.n294 30.8338
R3666 dvdd.n409 dvdd.n301 30.8338
R3667 dvdd.n562 dvdd.n301 30.8338
R3668 dvdd.n411 dvdd.n306 30.8338
R3669 dvdd.n556 dvdd.n306 30.8338
R3670 dvdd.n413 dvdd.n311 30.8338
R3671 dvdd.n550 dvdd.n311 30.8338
R3672 dvdd.n546 dvdd.n415 30.8338
R3673 dvdd.n422 dvdd.n415 30.8338
R3674 dvdd.n472 dvdd.n469 30.8338
R3675 dvdd.n477 dvdd.n472 30.8338
R3676 dvdd.n474 dvdd.n473 30.8338
R3677 dvdd.n477 dvdd.n473 30.8338
R3678 dvdd.n229 dvdd.n228 30.4946
R3679 dvdd.n183 dvdd.t213 29.5505
R3680 dvdd.n183 dvdd.t37 29.5505
R3681 dvdd.n239 dvdd.n178 29.3652
R3682 dvdd.n203 dvdd.n193 28.9887
R3683 dvdd.n201 dvdd.n200 28.6123
R3684 dvdd.n248 dvdd.n174 28.6123
R3685 dvdd.n288 dvdd.t42 28.5655
R3686 dvdd.n288 dvdd.t119 28.5655
R3687 dvdd.n209 dvdd.n208 27.4829
R3688 dvdd.n383 dvdd.n382 27.4147
R3689 dvdd.n383 dvdd.n339 27.4147
R3690 dvdd.n399 dvdd.n339 27.4147
R3691 dvdd.n400 dvdd.n399 27.4147
R3692 dvdd.n401 dvdd.n400 27.4147
R3693 dvdd.n401 dvdd.n290 27.4147
R3694 dvdd.n570 dvdd.n291 27.4147
R3695 dvdd.n560 dvdd.n291 27.4147
R3696 dvdd.n560 dvdd.n559 27.4147
R3697 dvdd.n559 dvdd.n558 27.4147
R3698 dvdd.n558 dvdd.n304 27.4147
R3699 dvdd.n548 dvdd.n304 27.4147
R3700 dvdd.n263 dvdd.n170 26.7299
R3701 dvdd.n479 dvdd.n478 26.4291
R3702 dvdd.n476 dvdd.n475 26.4291
R3703 dvdd.n177 dvdd.t127 26.3844
R3704 dvdd.n173 dvdd.t133 26.3844
R3705 dvdd.n172 dvdd.t123 26.3844
R3706 dvdd.n168 dvdd.t129 26.3844
R3707 dvdd.n168 dvdd.t247 26.3844
R3708 dvdd.n261 dvdd.t245 26.3844
R3709 dvdd.n261 dvdd.t249 26.3844
R3710 dvdd.n215 dvdd.n214 25.977
R3711 dvdd.n263 dvdd.n262 25.977
R3712 dvdd.n481 dvdd.n480 25.7522
R3713 dvdd.t250 dvdd.t9 25.5993
R3714 dvdd.n252 dvdd.n174 24.8476
R3715 dvdd.n256 dvdd.n169 24.8476
R3716 dvdd.n262 dvdd.n169 24.8476
R3717 dvdd.n511 dvdd.n510 24.0701
R3718 dvdd.n510 dvdd.n509 24.0701
R3719 dvdd.n571 dvdd.n570 23.8871
R3720 dvdd.n248 dvdd.n247 23.7181
R3721 dvdd.t108 dvdd.t212 23.5428
R3722 dvdd.n382 dvdd.n381 23.3832
R3723 dvdd.n200 dvdd.n196 23.3417
R3724 dvdd.n244 dvdd.n178 23.3417
R3725 dvdd.t134 dvdd.t75 19.9107
R3726 dvdd.n256 dvdd.n255 18.824
R3727 dvdd.n591 dvdd.n587 18.5005
R3728 dvdd.n592 dvdd.n591 18.5005
R3729 dvdd.n609 dvdd.n608 18.5005
R3730 dvdd.n610 dvdd.n609 18.5005
R3731 dvdd.n603 dvdd.n600 18.5005
R3732 dvdd.n589 dvdd.n588 18.5005
R3733 dvdd.n456 dvdd.n455 18.5005
R3734 dvdd.n455 dvdd.n444 18.5005
R3735 dvdd.n459 dvdd.n458 18.5005
R3736 dvdd.n458 dvdd.n445 18.5005
R3737 dvdd.n524 dvdd.n523 18.5005
R3738 dvdd.n525 dvdd.n524 18.5005
R3739 dvdd.n519 dvdd.n492 18.5005
R3740 dvdd.n519 dvdd.n518 18.5005
R3741 dvdd.n449 dvdd.n448 18.5005
R3742 dvdd dvdd.t128 17.0664
R3743 dvdd.n255 dvdd.n254 16.1887
R3744 dvdd.n285 dvdd.n167 15.4358
R3745 dvdd.n506 dvdd.n496 15.4172
R3746 dvdd.n507 dvdd.n506 15.4172
R3747 dvdd.n499 dvdd.n497 15.4172
R3748 dvdd.n516 dvdd.n515 15.4172
R3749 dvdd.n517 dvdd.n516 15.4172
R3750 dvdd.n196 dvdd.n167 14.6829
R3751 dvdd.t287 dvdd.t320 14.6159
R3752 dvdd.n593 dvdd.n581 12.7398
R3753 dvdd.n613 dvdd.n582 12.7398
R3754 dvdd.n450 dvdd.n440 12.5612
R3755 dvdd.n105 dvdd.n97 11.8036
R3756 dvdd.n117 dvdd.n116 11.8036
R3757 dvdd.n163 dvdd.n162 11.6875
R3758 dvdd.n262 dvdd.n260 10.3029
R3759 dvdd.t169 dvdd.t219 10.0458
R3760 dvdd.t124 dvdd.t164 9.95559
R3761 dvdd.n247 dvdd.n246 9.78874
R3762 dvdd.n601 dvdd.n582 9.58533
R3763 dvdd.n614 dvdd.n581 9.52467
R3764 dvdd.n532 dvdd.n441 9.45097
R3765 dvdd.n464 dvdd.n441 9.45097
R3766 dvdd.n522 dvdd.n464 9.45097
R3767 dvdd.n522 dvdd.n521 9.45097
R3768 dvdd.n217 dvdd.n216 9.41227
R3769 dvdd.n279 dvdd.n170 9.41227
R3770 dvdd.n279 dvdd.n278 9.3005
R3771 dvdd.n264 dvdd.n263 9.3005
R3772 dvdd.n286 dvdd.n285 9.3005
R3773 dvdd.n197 dvdd.n167 9.3005
R3774 dvdd.n198 dvdd.n196 9.3005
R3775 dvdd.n200 dvdd.n199 9.3005
R3776 dvdd.n201 dvdd.n194 9.3005
R3777 dvdd.n204 dvdd.n203 9.3005
R3778 dvdd.n205 dvdd.n193 9.3005
R3779 dvdd.n208 dvdd.n206 9.3005
R3780 dvdd.n209 dvdd.n191 9.3005
R3781 dvdd.n211 dvdd.n210 9.3005
R3782 dvdd.n212 dvdd.n190 9.3005
R3783 dvdd.n214 dvdd.n213 9.3005
R3784 dvdd.n217 dvdd.n189 9.3005
R3785 dvdd.n219 dvdd.n218 9.3005
R3786 dvdd.n221 dvdd.n220 9.3005
R3787 dvdd.n223 dvdd.n185 9.3005
R3788 dvdd.n225 dvdd.n224 9.3005
R3789 dvdd.n226 dvdd.n184 9.3005
R3790 dvdd.n228 dvdd.n227 9.3005
R3791 dvdd.n230 dvdd.n182 9.3005
R3792 dvdd.n233 dvdd.n232 9.3005
R3793 dvdd.n235 dvdd.n234 9.3005
R3794 dvdd.n237 dvdd.n179 9.3005
R3795 dvdd.n241 dvdd.n240 9.3005
R3796 dvdd.n242 dvdd.n178 9.3005
R3797 dvdd.n244 dvdd.n243 9.3005
R3798 dvdd.n245 dvdd.n175 9.3005
R3799 dvdd.n249 dvdd.n248 9.3005
R3800 dvdd.n250 dvdd.n174 9.3005
R3801 dvdd.n252 dvdd.n251 9.3005
R3802 dvdd.n253 dvdd.n171 9.3005
R3803 dvdd.n257 dvdd.n256 9.3005
R3804 dvdd.n258 dvdd.n169 9.3005
R3805 dvdd.t160 dvdd.n282 9.12162
R3806 dvdd.t248 dvdd.t0 8.53343
R3807 dvdd.n604 dvdd.t176 7.19008
R3808 dvdd.t67 dvdd.t110 7.11128
R3809 dvdd.n164 dvdd.n143 6.95702
R3810 dvdd.n512 dvdd.n489 6.69957
R3811 dvdd.n284 dvdd 5.938
R3812 dvdd.n513 dvdd.n512 5.74256
R3813 dvdd.t171 dvdd.t217 5.68912
R3814 dvdd.n230 dvdd.n229 5.64756
R3815 dvdd.n479 dvdd.n471 5.32439
R3816 dvdd.n533 dvdd.n440 4.96499
R3817 dvdd.n475 dvdd 4.94493
R3818 dvdd.n470 dvdd 4.91498
R3819 dvdd.n221 dvdd.n188 4.89462
R3820 dvdd.n102 dvdd.n101 4.74409
R3821 dvdd.t96 dvdd.n102 4.74409
R3822 dvdd.n104 dvdd.n103 4.74409
R3823 dvdd.n103 dvdd.t96 4.74409
R3824 dvdd.n112 dvdd.n110 4.74409
R3825 dvdd.t148 dvdd.n112 4.74409
R3826 dvdd.n111 dvdd.n109 4.74409
R3827 dvdd.t148 dvdd.n111 4.74409
R3828 dvdd.n164 dvdd.n163 4.73093
R3829 dvdd.n262 dvdd.n259 4.6255
R3830 dvdd.n500 dvdd.t335 4.61562
R3831 dvdd.n546 dvdd.n545 4.58635
R3832 dvdd.n533 dvdd.n532 4.48648
R3833 dvdd.n113 dvdd.n108 4.4805
R3834 dvdd.n98 dvdd.n96 4.3205
R3835 dvdd.t141 dvdd.t242 4.26697
R3836 dvdd.n236 dvdd.n235 4.14168
R3837 dvdd.n484 dvdd.n483 3.72349
R3838 dvdd.n118 dvdd.n108 3.64533
R3839 dvdd.n106 dvdd.n96 3.64377
R3840 dvdd.n571 dvdd.n290 3.52806
R3841 dvdd.n614 dvdd.n613 3.21567
R3842 dvdd.n489 dvdd.n488 2.7605
R3843 dvdd.n521 dvdd.n489 2.7519
R3844 dvdd.n240 dvdd.n238 2.63579
R3845 dvdd.n246 dvdd.n245 2.63579
R3846 dvdd.n105 dvdd.n104 2.55599
R3847 dvdd.n117 dvdd.n109 2.55599
R3848 dvdd.n480 dvdd.n470 2.28621
R3849 dvdd.n203 dvdd.n201 1.88285
R3850 dvdd.n277 dvdd.n276 1.8605
R3851 dvdd.n481 dvdd.n469 1.81103
R3852 dvdd.t325 dvdd.t327 1.42266
R3853 dvdd.n287 dvdd.n286 1.34131
R3854 dvdd.n254 dvdd.n253 1.12991
R3855 dvdd.n482 dvdd.n481 1.03383
R3856 dvdd.n165 dvdd.n164 1.01717
R3857 dvdd.n534 dvdd.n533 1.01588
R3858 dvdd.n82 dvdd 0.88709
R3859 dvdd dvdd.n277 0.877536
R3860 dvdd.n216 dvdd.n215 0.753441
R3861 dvdd.n222 dvdd.n221 0.753441
R3862 dvdd.n231 dvdd.n230 0.753441
R3863 dvdd.n240 dvdd.n239 0.753441
R3864 dvdd.n277 dvdd.n266 0.7505
R3865 dvdd.n543 dvdd.n535 0.687587
R3866 dvdd.n136 dvdd.n135 0.536822
R3867 dvdd.n578 dvdd.n287 0.53452
R3868 dvdd.n135 dvdd.n134 0.462454
R3869 dvdd.n287 dvdd 0.442652
R3870 dvdd.n615 dvdd.n614 0.423478
R3871 dvdd.n580 dvdd.n139 0.420507
R3872 dvdd.n514 dvdd.n513 0.419192
R3873 dvdd.n535 dvdd.n437 0.409354
R3874 dvdd.n579 dvdd.n140 0.407877
R3875 dvdd.n579 dvdd.n578 0.401019
R3876 dvdd.n487 dvdd.n467 0.40101
R3877 dvdd.n466 dvdd.n465 0.397184
R3878 dvdd.n439 dvdd.n438 0.392082
R3879 dvdd.n137 dvdd.n0 0.386761
R3880 dvdd.n616 dvdd.n138 0.386061
R3881 dvdd.n208 dvdd.n193 0.376971
R3882 dvdd.n235 dvdd.n181 0.376971
R3883 dvdd.n576 dvdd.n575 0.362045
R3884 dvdd.n136 dvdd.n1 0.359532
R3885 dvdd.n134 dvdd.t118 0.352122
R3886 dvdd.n486 dvdd.n485 0.349285
R3887 dvdd.n486 dvdd.n468 0.316676
R3888 dvdd.n487 dvdd.n486 0.29878
R3889 dvdd.n135 dvdd.n133 0.294897
R3890 dvdd.n480 dvdd.n479 0.283686
R3891 dvdd.n134 dvdd.t349 0.240872
R3892 dvdd.n572 dvdd.n571 0.226338
R3893 dvdd.n276 dvdd.n275 0.210336
R3894 dvdd.n433 dvdd.n432 0.209789
R3895 dvdd.n466 dvdd.n439 0.207511
R3896 dvdd.n544 dvdd.n543 0.202537
R3897 dvdd.n543 dvdd.n542 0.197568
R3898 dvdd.n535 dvdd.n534 0.194944
R3899 dvdd.n427 dvdd.n426 0.18972
R3900 dvdd.n82 dvdd.n81 0.188
R3901 dvdd.n84 dvdd.n79 0.188
R3902 dvdd.n86 dvdd.n73 0.188
R3903 dvdd.n88 dvdd.n67 0.188
R3904 dvdd.n90 dvdd.n61 0.188
R3905 dvdd.n92 dvdd.n55 0.188
R3906 dvdd.n94 dvdd.n49 0.188
R3907 dvdd.n120 dvdd.n43 0.188
R3908 dvdd.n122 dvdd.n37 0.188
R3909 dvdd.n124 dvdd.n31 0.188
R3910 dvdd.n126 dvdd.n25 0.188
R3911 dvdd.n128 dvdd.n19 0.188
R3912 dvdd.n130 dvdd.n13 0.188
R3913 dvdd.n132 dvdd.n7 0.188
R3914 dvdd.n133 dvdd.n4 0.188
R3915 dvdd.n131 dvdd.n10 0.188
R3916 dvdd.n129 dvdd.n16 0.188
R3917 dvdd.n127 dvdd.n22 0.188
R3918 dvdd.n125 dvdd.n28 0.188
R3919 dvdd.n123 dvdd.n34 0.188
R3920 dvdd.n121 dvdd.n40 0.188
R3921 dvdd.n95 dvdd.n46 0.188
R3922 dvdd.n93 dvdd.n52 0.188
R3923 dvdd.n91 dvdd.n58 0.188
R3924 dvdd.n89 dvdd.n64 0.188
R3925 dvdd.n87 dvdd.n70 0.188
R3926 dvdd.n85 dvdd.n76 0.188
R3927 dvdd.n83 dvdd.n80 0.188
R3928 dvdd.n429 dvdd.n428 0.183413
R3929 dvdd.n431 dvdd.n430 0.181119
R3930 dvdd.n488 dvdd 0.165183
R3931 dvdd.n540 dvdd.n539 0.158073
R3932 dvdd.n538 dvdd.n537 0.157259
R3933 dvdd.n166 dvdd.n165 0.155583
R3934 dvdd.n264 dvdd.n259 0.154565
R3935 dvdd.n536 dvdd.n289 0.153187
R3936 dvdd.n542 dvdd.n541 0.153187
R3937 dvdd.n574 dvdd.n573 0.151151
R3938 dvdd.n575 dvdd.n574 0.148301
R3939 dvdd.n430 dvdd.n429 0.134674
R3940 dvdd dvdd.n166 0.129649
R3941 dvdd.n428 dvdd.n427 0.126647
R3942 dvdd.n426 dvdd.n425 0.121486
R3943 dvdd.n545 dvdd.n434 0.121486
R3944 dvdd.n432 dvdd.n431 0.116326
R3945 dvdd.n580 dvdd.n579 0.111459
R3946 dvdd.n119 dvdd.n118 0.105151
R3947 dvdd.n107 dvdd.n106 0.105151
R3948 dvdd.n259 dvdd 0.103283
R3949 dvdd.n198 dvdd.n197 0.103064
R3950 dvdd.n199 dvdd.n198 0.103064
R3951 dvdd.n199 dvdd.n194 0.103064
R3952 dvdd.n204 dvdd.n194 0.103064
R3953 dvdd.n205 dvdd.n204 0.103064
R3954 dvdd.n206 dvdd.n205 0.103064
R3955 dvdd.n206 dvdd.n191 0.103064
R3956 dvdd.n211 dvdd.n191 0.103064
R3957 dvdd.n212 dvdd.n211 0.103064
R3958 dvdd.n213 dvdd.n212 0.103064
R3959 dvdd.n213 dvdd.n189 0.103064
R3960 dvdd.n219 dvdd.n189 0.103064
R3961 dvdd.n220 dvdd.n219 0.103064
R3962 dvdd.n220 dvdd.n185 0.103064
R3963 dvdd.n225 dvdd.n185 0.103064
R3964 dvdd.n226 dvdd.n225 0.103064
R3965 dvdd.n227 dvdd.n226 0.103064
R3966 dvdd.n227 dvdd.n182 0.103064
R3967 dvdd.n233 dvdd.n182 0.103064
R3968 dvdd.n234 dvdd.n233 0.103064
R3969 dvdd.n234 dvdd.n179 0.103064
R3970 dvdd.n241 dvdd.n179 0.103064
R3971 dvdd.n243 dvdd.n242 0.103064
R3972 dvdd.n243 dvdd.n175 0.103064
R3973 dvdd.n249 dvdd.n175 0.103064
R3974 dvdd.n250 dvdd.n249 0.103064
R3975 dvdd.n251 dvdd.n250 0.103064
R3976 dvdd.n251 dvdd.n171 0.103064
R3977 dvdd.n257 dvdd.n171 0.103064
R3978 dvdd.n534 dvdd.n439 0.0977222
R3979 dvdd.n434 dvdd.n433 0.0974037
R3980 dvdd.n266 dvdd.n265 0.0907869
R3981 dvdd.n137 dvdd.n136 0.0905685
R3982 dvdd.n577 dvdd.n576 0.0820092
R3983 dvdd.n537 dvdd.n536 0.0693111
R3984 dvdd.n541 dvdd.n540 0.0664609
R3985 dvdd.n539 dvdd.n538 0.0660537
R3986 dvdd.n545 dvdd.n544 0.0635734
R3987 dvdd.n615 dvdd.n580 0.0611164
R3988 dvdd.n265 dvdd 0.0568119
R3989 dvdd.n286 dvdd 0.0517821
R3990 dvdd.n197 dvdd 0.0517821
R3991 dvdd dvdd.n241 0.0517821
R3992 dvdd.n242 dvdd 0.0517821
R3993 dvdd dvdd.n257 0.0517821
R3994 dvdd.n258 dvdd 0.0517821
R3995 dvdd dvdd.n258 0.0517821
R3996 dvdd dvdd.n264 0.0517821
R3997 dvdd.n278 dvdd 0.0517821
R3998 dvdd.n278 dvdd 0.0517821
R3999 dvdd.n573 dvdd.n572 0.0505814
R4000 dvdd.n485 dvdd.n484 0.048322
R4001 dvdd.n483 dvdd 0.0436596
R4002 dvdd.n578 dvdd.n577 0.0425507
R4003 dvdd.n84 dvdd.n83 0.0386466
R4004 dvdd.n86 dvdd.n85 0.0386466
R4005 dvdd.n88 dvdd.n87 0.0386466
R4006 dvdd.n90 dvdd.n89 0.0386466
R4007 dvdd.n92 dvdd.n91 0.0386466
R4008 dvdd.n94 dvdd.n93 0.0386466
R4009 dvdd.n122 dvdd.n121 0.0386466
R4010 dvdd.n124 dvdd.n123 0.0386466
R4011 dvdd.n126 dvdd.n125 0.0386466
R4012 dvdd.n128 dvdd.n127 0.0386466
R4013 dvdd.n130 dvdd.n129 0.0386466
R4014 dvdd.n132 dvdd.n131 0.0386466
R4015 dvdd dvdd.n137 0.0316644
R4016 dvdd dvdd.n466 0.0296005
R4017 dvdd.n107 dvdd.n95 0.0295948
R4018 dvdd dvdd.n616 0.0237877
R4019 dvdd.n616 dvdd.n615 0.0234452
R4020 dvdd.n488 dvdd.n487 0.0196799
R4021 dvdd.n572 dvdd.n289 0.0180081
R4022 dvdd.n106 dvdd.n105 0.0173379
R4023 dvdd.n118 dvdd.n117 0.0173379
R4024 dvdd.n120 dvdd.n119 0.00631897
R4025 dvdd.n483 dvdd.n482 0.0041645
R4026 dvdd.n83 dvdd.n82 0.00373276
R4027 dvdd.n85 dvdd.n84 0.00373276
R4028 dvdd.n87 dvdd.n86 0.00373276
R4029 dvdd.n89 dvdd.n88 0.00373276
R4030 dvdd.n91 dvdd.n90 0.00373276
R4031 dvdd.n93 dvdd.n92 0.00373276
R4032 dvdd.n95 dvdd.n94 0.00373276
R4033 dvdd.n119 dvdd.n107 0.00373276
R4034 dvdd.n121 dvdd.n120 0.00373276
R4035 dvdd.n123 dvdd.n122 0.00373276
R4036 dvdd.n125 dvdd.n124 0.00373276
R4037 dvdd.n127 dvdd.n126 0.00373276
R4038 dvdd.n129 dvdd.n128 0.00373276
R4039 dvdd.n131 dvdd.n130 0.00373276
R4040 dvdd.n133 dvdd.n132 0.00373276
R4041 dvdd.n482 dvdd 0.00131433
R4042 a_35262_n291454.t24 a_35262_n291454.t29 353.467
R4043 a_35262_n291454.t15 a_35262_n291454.t23 353.467
R4044 a_35262_n291454.t12 a_35262_n291454.t18 353.467
R4045 a_35262_n291454.t21 a_35262_n291454.t27 353.467
R4046 a_35262_n291454.t7 a_35262_n291454.t11 353.467
R4047 a_35262_n291454.t17 a_35262_n291454.t25 353.467
R4048 a_35262_n291454.t26 a_35262_n291454.t6 353.467
R4049 a_35262_n291454.t10 a_35262_n291454.t16 353.467
R4050 a_35262_n291454.n18 a_35262_n291454.n0 299.851
R4051 a_35262_n291454.n19 a_35262_n291454.n18 299.414
R4052 a_35262_n291454.n2 a_35262_n291454.t24 232.382
R4053 a_35262_n291454.n5 a_35262_n291454.t10 232.382
R4054 a_35262_n291454.n17 a_35262_n291454.n1 197.161
R4055 a_35262_n291454.n12 a_35262_n291454.t8 185.79
R4056 a_35262_n291454.n9 a_35262_n291454.t19 185.79
R4057 a_35262_n291454.n2 a_35262_n291454.t15 162.274
R4058 a_35262_n291454.n3 a_35262_n291454.t12 162.274
R4059 a_35262_n291454.n4 a_35262_n291454.t21 162.274
R4060 a_35262_n291454.n7 a_35262_n291454.t7 162.274
R4061 a_35262_n291454.n6 a_35262_n291454.t17 162.274
R4062 a_35262_n291454.n5 a_35262_n291454.t26 162.274
R4063 a_35262_n291454.n12 a_35262_n291454.t22 115.68
R4064 a_35262_n291454.n13 a_35262_n291454.t14 115.68
R4065 a_35262_n291454.n14 a_35262_n291454.t28 115.68
R4066 a_35262_n291454.n11 a_35262_n291454.t20 115.68
R4067 a_35262_n291454.n10 a_35262_n291454.t9 115.68
R4068 a_35262_n291454.n9 a_35262_n291454.t13 115.68
R4069 a_35262_n291454.n10 a_35262_n291454.n9 70.1096
R4070 a_35262_n291454.n11 a_35262_n291454.n10 70.1096
R4071 a_35262_n291454.n14 a_35262_n291454.n13 70.1096
R4072 a_35262_n291454.n13 a_35262_n291454.n12 70.1096
R4073 a_35262_n291454.n3 a_35262_n291454.n2 70.1096
R4074 a_35262_n291454.n4 a_35262_n291454.n3 70.1096
R4075 a_35262_n291454.n7 a_35262_n291454.n6 70.1096
R4076 a_35262_n291454.n6 a_35262_n291454.n5 70.1096
R4077 a_35262_n291454.n0 a_35262_n291454.t2 46.4362
R4078 a_35262_n291454.n0 a_35262_n291454.t4 46.4362
R4079 a_35262_n291454.n19 a_35262_n291454.t3 46.4362
R4080 a_35262_n291454.t5 a_35262_n291454.n19 46.4362
R4081 a_35262_n291454.n1 a_35262_n291454.t1 39.6005
R4082 a_35262_n291454.n1 a_35262_n291454.t0 39.6005
R4083 a_35262_n291454.n15 a_35262_n291454.n11 35.055
R4084 a_35262_n291454.n15 a_35262_n291454.n14 35.055
R4085 a_35262_n291454.n8 a_35262_n291454.n4 35.055
R4086 a_35262_n291454.n8 a_35262_n291454.n7 35.055
R4087 a_35262_n291454.n16 a_35262_n291454.n15 17.6874
R4088 a_35262_n291454.n16 a_35262_n291454.n8 17.6491
R4089 a_35262_n291454.n17 a_35262_n291454.n16 2.43319
R4090 a_35262_n291454.n18 a_35262_n291454.n17 0.572285
R4091 x2.Td_Sd.t6 x2.Td_Sd.t7 1548.83
R4092 x2.Td_Sd.t7 x2.Td_Sd.n1 355.707
R4093 x2.Td_Sd.n13 x2.Td_Sd.t1 346.822
R4094 x2.Td_Sd.n11 x2.Td_Sd.t5 346.644
R4095 x2.Td_Sd.n11 x2.Td_Sd.t0 345.853
R4096 x2.Td_Sd.n13 x2.Td_Sd.t2 345.849
R4097 x2.Td_Sd.n0 x2.Td_Sd.t16 295.091
R4098 x2.Td_Sd.n8 x2.Td_Sd.t8 272.087
R4099 x2.Td_Sd.n6 x2.Td_Sd.t12 250.909
R4100 x2.Td_Sd.n4 x2.Td_Sd.t10 241
R4101 x2.Td_Sd.n14 x2.Td_Sd.t4 236.911
R4102 x2.Td_Sd.n12 x2.Td_Sd.t3 236.799
R4103 x2.Td_Sd.n0 x2.Td_Sd.t11 236.18
R4104 x2.Td_Sd.n1 x2.Td_Sd.t13 227.27
R4105 x2.Td_Sd.n2 x2.Td_Sd.t6 204.88
R4106 x2.Td_Sd.n6 x2.Td_Sd.t17 199.227
R4107 x2.Td_Sd.n8 x2.Td_Sd.t14 184.476
R4108 x2.Td_Sd.n2 x2.Td_Sd.t9 184.369
R4109 x2.Td_Sd.n4 x2.Td_Sd.t15 176.588
R4110 x2.Td_Sd.n9 x2.Td_Sd.n8 176.243
R4111 x2.Td_Sd.n3 x2.Td_Sd.n0 169.823
R4112 x2.Td_Sd.n3 x2.Td_Sd.n2 162.852
R4113 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtp_1_0.CLK x2.Td_Sd.n4 156.542
R4114 x2.Td_Sd.n7 x2.Td_Sd.n6 152
R4115 x2.Td_Sd.n7 x2.delayPulse_digital_0/sky130_fd_sc_ls__xor2_1_0.B 18.824
R4116 x2.Td_Sd.n9 x2.delayPulse_digital_0/sky130_fd_sc_ls__xor2_1_0.B 18.6187
R4117 x2.Td_Sd.n5 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtp_1_0.CLK 13.7738
R4118 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.RESET_B x2.Td_Sd.n1 159.315
R4119 x2.Td_Sd.n12 x2.Td_Sd.n10 12.4112
R4120 x2.Td_Sd.n10 x2.Td_Sd.n9 10.5303
R4121 x2.Td_Sd.n10 x2.Td_Sd.n5 6.2147
R4122 x2.delayPulse_digital_0/sky130_fd_sc_ls__xor2_1_0.B x2.Td_Sd.n7 4.84898
R4123 x2.Td_Sd.n14 x2.Td_Sd.n13 0.91089
R4124 x2.Td_Sd.n12 x2.Td_Sd.n11 0.745991
R4125 x2.Td_Sd.n14 x2.Td_Sd.n12 0.563933
R4126 x2.Td_Sd.n5 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.RESET_B 6.46049
R4127 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.RESET_B x2.Td_Sd.n3 3.32775
R4128 a_25883_n288267.n2 a_25883_n288267.t3 341.05
R4129 a_25883_n288267.t1 a_25883_n288267.n2 340.209
R4130 a_25883_n288267.n2 a_25883_n288267.t2 231.944
R4131 a_25883_n288267.n8 a_25883_n288267.t4 190.986
R4132 a_25883_n288267.t4 a_25883_n288267.n7 190.986
R4133 a_25883_n288267.n6 a_25883_n288267.t9 190.986
R4134 a_25883_n288267.t9 a_25883_n288267.n5 190.986
R4135 a_25883_n288267.t5 a_25883_n288267.n5 190.954
R4136 a_25883_n288267.n6 a_25883_n288267.t5 190.954
R4137 a_25883_n288267.n7 a_25883_n288267.t6 190.954
R4138 a_25883_n288267.n8 a_25883_n288267.t6 190.954
R4139 a_25883_n288267.n4 a_25883_n288267.t7 170.1
R4140 a_25883_n288267.t7 a_25883_n288267.n3 170.1
R4141 a_25883_n288267.t8 a_25883_n288267.n3 170.069
R4142 a_25883_n288267.n4 a_25883_n288267.t8 170.069
R4143 a_25883_n288267.n0 a_25883_n288267.n5 67.7619
R4144 a_25883_n288267.n1 a_25883_n288267.n3 67.7467
R4145 a_25883_n288267.n1 a_25883_n288267.n4 66.9702
R4146 a_25883_n288267.n0 a_25883_n288267.n6 66.9021
R4147 a_25883_n288267.n7 a_25883_n288267.n0 66.9021
R4148 a_25883_n288267.n0 a_25883_n288267.n8 66.9021
R4149 a_25883_n288267.n2 a_25883_n288267.t0 8.29364
R4150 a_25883_n288267.n2 a_25883_n288267.n1 2.76399
R4151 a_25883_n288267.n1 a_25883_n288267.n0 2.41607
R4152 a_36398_n287783.n0 a_36398_n287783.t6 157.31
R4153 a_36398_n287783.n0 a_36398_n287783.t7 157.31
R4154 a_36398_n287783.n0 a_36398_n287783.t4 119.243
R4155 a_36398_n287783.n0 a_36398_n287783.t5 119.243
R4156 a_36398_n287783.n2 a_36398_n287783.n1 86.5831
R4157 a_36398_n287783.n1 a_36398_n287783.t1 85.3779
R4158 a_36398_n287783.n1 a_36398_n287783.t3 85.227
R4159 a_36398_n287783.t0 a_36398_n287783.n2 11.0785
R4160 a_36398_n287783.n2 a_36398_n287783.t2 11.0785
R4161 a_36398_n287783.n1 a_36398_n287783.n0 1.97928
R4162 a_37002_n287783.n0 a_37002_n287783.t7 159.1
R4163 a_37002_n287783.n0 a_37002_n287783.t5 157.478
R4164 a_37002_n287783.n0 a_37002_n287783.t6 119.55
R4165 a_37002_n287783.n0 a_37002_n287783.t4 119.531
R4166 a_37002_n287783.n2 a_37002_n287783.n1 86.5435
R4167 a_37002_n287783.n1 a_37002_n287783.t0 85.3657
R4168 a_37002_n287783.n1 a_37002_n287783.t1 85.2346
R4169 a_37002_n287783.n2 a_37002_n287783.t3 11.0785
R4170 a_37002_n287783.t2 a_37002_n287783.n2 11.0785
R4171 a_37002_n287783.n1 a_37002_n287783.n0 2.06116
R4172 a_32918_n290853.n2 a_32918_n290853.t1 341.137
R4173 a_32918_n290853.t2 a_32918_n290853.n2 340.207
R4174 a_32918_n290853.n2 a_32918_n290853.t0 231.925
R4175 a_32918_n290853.n6 a_32918_n290853.t6 190.986
R4176 a_32918_n290853.t6 a_32918_n290853.n5 190.986
R4177 a_32918_n290853.n4 a_32918_n290853.t8 190.986
R4178 a_32918_n290853.t8 a_32918_n290853.n3 190.986
R4179 a_32918_n290853.t5 a_32918_n290853.n3 190.954
R4180 a_32918_n290853.n4 a_32918_n290853.t5 190.954
R4181 a_32918_n290853.n5 a_32918_n290853.t3 190.954
R4182 a_32918_n290853.n6 a_32918_n290853.t3 190.954
R4183 a_32918_n290853.n8 a_32918_n290853.t4 170.1
R4184 a_32918_n290853.t4 a_32918_n290853.n7 170.1
R4185 a_32918_n290853.t7 a_32918_n290853.n7 170.069
R4186 a_32918_n290853.n8 a_32918_n290853.t7 170.069
R4187 a_32918_n290853.n0 a_32918_n290853.n3 67.7868
R4188 a_32918_n290853.n1 a_32918_n290853.n7 67.6654
R4189 a_32918_n290853.n0 a_32918_n290853.n4 66.9439
R4190 a_32918_n290853.n5 a_32918_n290853.n0 66.9439
R4191 a_32918_n290853.n1 a_32918_n290853.n6 66.9439
R4192 a_32918_n290853.n1 a_32918_n290853.n8 66.9225
R4193 a_32918_n290853.n1 a_32918_n290853.n0 2.01708
R4194 a_32918_n290853.n2 a_32918_n290853.n1 1.96404
R4195 x2.Td_L.t14 x2.Td_L.t10 803.333
R4196 x2.Td_L.t10 x2.Td_L.t11 484.947
R4197 x2.Td_L.n15 x2.Td_L.n13 300.317
R4198 x2.Td_L.n15 x2.Td_L.n14 299.408
R4199 x2.Td_L.n7 x2.Td_L.t7 260.281
R4200 x2.Td_L x2.Td_L.n12 197.181
R4201 x2.Td_L.t8 x2.Td_L.n9 190.986
R4202 x2.Td_L.n6 x2.Td_L.t12 190.986
R4203 x2.Td_L.t12 x2.Td_L.n5 190.986
R4204 x2.Td_L.t6 x2.Td_L.n5 190.954
R4205 x2.Td_L.n6 x2.Td_L.t6 190.954
R4206 x2.Td_L.n9 x2.Td_L.t13 190.954
R4207 x2.Td_L.n7 x2.Td_L.t14 173.228
R4208 x2.Td_L.n11 x2.Td_L.t15 170.1
R4209 x2.Td_L.t15 x2.Td_L.n10 170.1
R4210 x2.Td_L.t9 x2.Td_L.n10 170.069
R4211 x2.Td_L.n11 x2.Td_L.t9 170.069
R4212 x2.Td_L.n3 x2.Td_L.t8 190.969
R4213 x2.Td_L.n3 x2.Td_L.t13 190.969
R4214 x2.Td_L.n2 x2.Td_L.n3 66.3047
R4215 x2.Td_L.n8 x2.Td_L.n7 104.355
R4216 x2.Td_L.n4 x2.Td_L.n5 67.7404
R4217 x2.Td_L.n1 x2.Td_L.n10 67.6296
R4218 x2.Td_L.n4 x2.Td_L.n6 66.9082
R4219 x2.Td_L.n9 x2.Td_L.n4 66.9082
R4220 x2.Td_L.n1 x2.Td_L.n11 66.8868
R4221 x2.Td_L.n13 x2.Td_L.t2 46.4362
R4222 x2.Td_L.n13 x2.Td_L.t4 46.4362
R4223 x2.Td_L.n14 x2.Td_L.t3 46.4362
R4224 x2.Td_L.n14 x2.Td_L.t5 46.4362
R4225 x2.Td_L.n12 x2.Td_L.t1 39.6005
R4226 x2.Td_L.n12 x2.Td_L.t0 39.6005
R4227 x2.Td_L.n2 x2.Td_L.n8 37.5228
R4228 x2.Td_L x2.Td_L.n1 1.38176
R4229 x2.Td_L.n0 x2.Td_L.n4 1.09336
R4230 x2.Td_L.n1 x2.Td_L.n0 0.893357
R4231 x2.Td_L x2.Td_L.n15 0.891776
R4232 x2.Td_L.n0 x2.Td_L.n2 0.800888
R4233 x2.Td_L.n8 x2.Td_L 0.705087
R4234 a_4566_n291516.n0 a_4566_n291516.t2 227.352
R4235 a_4566_n291516.n1 a_4566_n291516.t3 196.169
R4236 a_4566_n291516.t0 a_4566_n291516.n1 23.6417
R4237 a_4566_n291516.n0 a_4566_n291516.t1 13.584
R4238 a_4566_n291516.n1 a_4566_n291516.n0 1.59969
R4239 x1.vbn.n5 x1.vbn.t6 264.832
R4240 x1.vbn.n0 x1.vbn.t0 230.387
R4241 x1.vbn.n6 x1.vbn.t7 72.4418
R4242 x1.vbn.n3 x1.vbn.t10 72.3203
R4243 x1.vbn.n2 x1.vbn.t5 72.3144
R4244 x1.vbn.n0 x1.vbn.t1 71.4758
R4245 x1.vbn.n2 x1.vbn.t4 70.7106
R4246 x1.vbn.n3 x1.vbn.t8 70.7033
R4247 x1.vbn.n6 x1.vbn.t9 70.6707
R4248 x1.vbn.n0 x1.vbn.t2 40.9588
R4249 x1.vbn.n5 x1.vbn.t3 23.5181
R4250 x1.vbn x1.vbn.n4 3.85926
R4251 x1.vbn.n4 x1.vbn.n2 2.92849
R4252 x1.vbn x1.vbn.n1 2.48447
R4253 x1.vbn.n1 x1.vbn.n5 2.22005
R4254 x1.vbn.n1 x1.vbn.n6 1.99442
R4255 x1.vbn.n4 x1.vbn.n3 1.88535
R4256 x1.vbn.n1 x1.vbn.n0 1.69839
R4257 a_5972_n290308.n0 a_5972_n290308.t4 228.429
R4258 a_5972_n290308.n0 a_5972_n290308.t0 41.8804
R4259 a_5972_n290308.n0 a_5972_n290308.t1 40.9588
R4260 a_5972_n290308.t2 a_5972_n290308.n1 23.5738
R4261 a_5972_n290308.n0 a_5972_n290308.t3 12.8438
R4262 a_5972_n290308.n1 a_5972_n290308.t5 12.8184
R4263 a_5972_n290308.n1 a_5972_n290308.n0 4.91266
R4264 avss.n214 avss.n200 325390
R4265 avss.n1047 avss.n1026 126229
R4266 avss.n1047 avss.n1027 120611
R4267 avss.n1231 avss.t13 113252
R4268 avss.n891 avss.n219 93411
R4269 avss.n1043 avss.n1027 93404.6
R4270 avss.n1043 avss.n1030 77113.4
R4271 avss.n1215 avss.t0 60898.5
R4272 avss.n1034 avss.n1026 54654.1
R4273 avss.t69 avss.n1231 42915.9
R4274 avss.n175 avss.n159 42361.3
R4275 avss.n552 avss.n505 40791.1
R4276 avss.n891 avss.n218 37112.5
R4277 avss.n1256 avss.n1255 33058.4
R4278 avss.n1034 avss.n1030 32711.6
R4279 avss.n1046 avss.n1028 29011.1
R4280 avss.n1082 avss.n161 25407.2
R4281 avss.n1086 avss.n161 25407.2
R4282 avss.n1086 avss.n162 25407.2
R4283 avss.n172 avss.n170 25407.2
R4284 avss.n174 avss.n172 25407.2
R4285 avss.n1073 avss.n170 25407.2
R4286 avss.n1073 avss.n174 25407.2
R4287 avss.n1046 avss.n1045 23251
R4288 avss.n1033 avss.n1028 22647.7
R4289 avss.n1243 avss.n25 21160.1
R4290 avss.n1254 avss.n25 21160.1
R4291 avss.n1243 avss.n26 21160.1
R4292 avss.n1254 avss.n26 21160.1
R4293 avss.n1045 avss.n1044 20409.5
R4294 avss.n148 avss.n143 16351
R4295 avss.n144 avss.n143 16351
R4296 avss.n148 avss.n146 16351
R4297 avss.n146 avss.n144 16351
R4298 avss.n920 avss.n893 16125.8
R4299 avss.n1072 avss.n1071 13403.5
R4300 avss.n775 avss.n768 13338.5
R4301 avss.n893 avss.n215 12361.9
R4302 avss.n890 avss.n889 11682.6
R4303 avss.n398 avss.n397 11392.7
R4304 avss.n500 avss.n499 10626
R4305 avss.n1090 avss.n1089 10436.2
R4306 avss.n892 avss.n891 10051.9
R4307 avss.n1071 avss.n175 9855.53
R4308 avss.n552 avss.n551 9608.16
R4309 avss.n1228 avss.n42 9322.74
R4310 avss.n1228 avss.n43 9322.74
R4311 avss.n1207 avss.n42 9322.74
R4312 avss.n1207 avss.n43 9322.74
R4313 avss.n601 avss.n501 9270.59
R4314 avss.n601 avss.n502 9270.59
R4315 avss.n595 avss.n502 9270.59
R4316 avss.n595 avss.n501 9270.59
R4317 avss.n550 avss.n507 9270.59
R4318 avss.n544 avss.n507 9270.59
R4319 avss.n550 avss.n508 9270.59
R4320 avss.n544 avss.n508 9270.59
R4321 avss.n553 avss.n552 9139.67
R4322 avss.n1159 avss.n75 9038.82
R4323 avss.n76 avss.n75 9038.82
R4324 avss.n1159 avss.n78 9038.82
R4325 avss.n78 avss.n76 9038.82
R4326 avss.n214 avss.n213 9007.72
R4327 avss.n659 avss.n658 8593.75
R4328 avss.n215 avss.n214 8503.42
R4329 avss.n20 avss.n6 8190.47
R4330 avss.n1044 avss.n1029 7497.54
R4331 avss.n505 avss.n217 7283.07
R4332 avss.n891 avss.n890 6982.95
R4333 avss.n893 avss.n892 5709.96
R4334 avss.n50 avss.n6 5683.2
R4335 avss.n775 avss.n159 5423.26
R4336 avss.n1148 avss.n82 5168.35
R4337 avss.n1149 avss.n82 5168.35
R4338 avss.n1235 avss.n38 5168.35
R4339 avss.n1236 avss.n38 5168.35
R4340 avss.n1079 avss.n163 5140.55
R4341 avss.n1091 avss.n1090 4970.28
R4342 avss.n811 dvss 4834.33
R4343 avss.n1090 avss.n136 4803
R4344 avss.n342 avss.n220 4692.56
R4345 avss.n1223 avss.n1222 4439.33
R4346 avss.n1062 avss.n181 4152.6
R4347 avss.n1062 avss.n182 4152.6
R4348 avss.n1258 avss.n14 4131.21
R4349 avss.n1258 avss.n23 4131.21
R4350 avss.n1257 avss.n14 4131.21
R4351 avss.n1257 avss.n23 4131.21
R4352 avss.n812 dvss 4092.31
R4353 avss.n1221 avss.n52 4025.74
R4354 dvss avss.n812 4018.54
R4355 avss.n1095 avss.n118 4018.37
R4356 avss.n551 avss.n506 3896.99
R4357 avss.n543 avss.n506 3896.99
R4358 avss.n602 avss.n601 3867.64
R4359 avss.n1033 avss.n1029 3860.74
R4360 avss.n1240 avss.n33 3760.38
R4361 avss.n1240 avss.n34 3760.38
R4362 avss.n1162 avss.n66 3760.38
R4363 avss.n70 avss.n66 3760.38
R4364 avss.n84 avss.n67 3760.38
R4365 avss.n84 avss.n83 3760.38
R4366 avss.n811 avss.n219 3686.18
R4367 avss.n217 avss.n215 3474.37
R4368 avss.n659 dvss 3413.97
R4369 avss.n477 avss.n220 3396.49
R4370 avss.n1211 avss.n1210 3115.28
R4371 avss.n1211 avss.n56 3115.28
R4372 avss.n1119 avss.n103 3115.28
R4373 avss.n1121 avss.n99 3115.28
R4374 avss.n1122 avss.n99 3115.28
R4375 avss.n1118 avss.n103 3115.28
R4376 avss.n61 avss.n56 3098.81
R4377 avss.n1210 avss.n61 3098.81
R4378 avss.n918 avss.n896 3075.76
R4379 avss.n918 avss.n895 3075.76
R4380 avss.n900 avss.n182 2953.91
R4381 avss.n905 avss.n181 2953.91
R4382 avss.n136 avss.n135 2634.65
R4383 avss.n1262 avss.n8 2575.21
R4384 avss.n1263 avss.n8 2575.21
R4385 avss.n1263 avss.n7 2575.21
R4386 avss.n1262 avss.n7 2575.21
R4387 avss.n1112 avss.n114 2575.21
R4388 avss.n1112 avss.n115 2575.21
R4389 avss.n1113 avss.n115 2575.21
R4390 avss.n1113 avss.n114 2575.21
R4391 avss.n1137 avss.n91 2575.21
R4392 avss.n1136 avss.n91 2575.21
R4393 avss.n1131 avss.n1130 2575.21
R4394 avss.n1132 avss.n1131 2575.21
R4395 avss.n928 avss.n197 2445.12
R4396 avss.n930 avss.n197 2445.12
R4397 avss.n935 avss.n188 2445.12
R4398 avss.n937 avss.n188 2445.12
R4399 avss.n923 avss.n207 2445.12
R4400 avss.n923 avss.n208 2445.12
R4401 avss.n776 avss.n774 2445.12
R4402 avss.n777 avss.n776 2445.12
R4403 avss.n157 avss.n137 2390.79
R4404 avss.n151 avss.n137 2390.79
R4405 avss.n157 avss.n138 2390.79
R4406 avss.n151 avss.n138 2390.79
R4407 avss.n540 avss.n512 2317.65
R4408 avss.n540 avss.n513 2317.65
R4409 avss.n804 avss.n734 2317.65
R4410 avss.n804 avss.n735 2317.65
R4411 avss.n1120 avss.n102 2216.26
R4412 avss.n102 avss.n98 2216.26
R4413 avss.n614 avss.n237 2127.34
R4414 avss.n628 avss.n237 2127.34
R4415 avss.n1216 avss.n53 2064.78
R4416 avss.n1216 avss.n54 2064.78
R4417 avss.n1219 avss.n54 2064.78
R4418 avss.n1219 avss.n53 2064.78
R4419 avss.n623 avss.n622 2041.29
R4420 avss.n227 avss.n221 2016.35
R4421 avss.n880 avss.n227 2016.35
R4422 avss.n888 avss.n224 2016.35
R4423 avss.n884 avss.n224 2016.35
R4424 avss.n808 avss.n656 2016.35
R4425 avss.n808 avss.n657 2016.35
R4426 avss.n816 avss.n656 2016.35
R4427 avss.n816 avss.n657 2016.35
R4428 avss.n892 avss.n216 1890.37
R4429 avss.n899 avss.n896 1877.07
R4430 avss.n903 avss.n895 1877.07
R4431 avss.n556 avss.n554 1863.9
R4432 avss.n592 avss.n556 1863.9
R4433 avss.n584 avss.n563 1863.9
R4434 avss.n584 avss.n564 1863.9
R4435 avss.n1125 avss.n92 1857.31
R4436 avss.n1125 avss.n95 1857.31
R4437 avss.n911 avss.n180 1836.58
R4438 avss.n1063 avss.n180 1836.58
R4439 avss.n624 avss.n604 1834.26
R4440 avss.n658 avss.n218 1797.26
R4441 avss.n1049 avss.n1024 1772.77
R4442 avss.n1069 avss.n177 1735.47
R4443 avss.n1069 avss.n178 1735.47
R4444 avss.n1065 avss.n178 1735.47
R4445 avss.n1065 avss.n177 1735.47
R4446 avss.n1048 avss.n1025 1653.19
R4447 avss.n1074 avss.n169 1650.89
R4448 avss.n1084 avss.n1083 1650.82
R4449 avss.n806 dvss 1628.88
R4450 avss.n1195 avss.n1191 1603.74
R4451 avss.n1194 avss.n1191 1603.74
R4452 avss.n1184 avss.n1182 1603.74
R4453 avss.n1185 avss.n1182 1603.74
R4454 avss.n134 avss.n129 1603.74
R4455 avss.n1099 avss.n1097 1603.74
R4456 avss.n1097 avss.n1094 1603.74
R4457 avss.n134 avss.n130 1603.74
R4458 avss.n809 avss.n806 1554.14
R4459 avss.n1071 avss.n1070 1539.06
R4460 avss.n615 avss.n238 1442.18
R4461 avss.n627 avss.n238 1442.18
R4462 avss.n1148 avss.n67 1407.97
R4463 avss.n1161 avss.n67 1407.97
R4464 avss.n1162 avss.n1161 1407.97
R4465 avss.n1163 avss.n1162 1407.97
R4466 avss.n1163 avss.n33 1407.97
R4467 avss.n1235 avss.n33 1407.97
R4468 avss.n1149 avss.n83 1407.97
R4469 avss.n83 avss.n71 1407.97
R4470 avss.n71 avss.n70 1407.97
R4471 avss.n70 avss.n69 1407.97
R4472 avss.n69 avss.n34 1407.97
R4473 avss.n1236 avss.n34 1407.97
R4474 avss.n928 avss.n201 1344.24
R4475 avss.n931 avss.n930 1344.24
R4476 avss.n935 avss.n192 1344.24
R4477 avss.n207 avss.n192 1344.24
R4478 avss.n937 avss.n189 1344.24
R4479 avss.n208 avss.n189 1344.24
R4480 avss.n784 avss.n756 1344.24
R4481 avss.n784 avss.n766 1344.24
R4482 avss.n774 avss.n766 1344.24
R4483 avss.n767 avss.n751 1344.24
R4484 avss.n769 avss.n767 1344.24
R4485 avss.n777 avss.n769 1344.24
R4486 avss.n50 avss.n49 1316.44
R4487 avss.n1042 avss.n1025 1305.96
R4488 avss.n542 avss.n505 1303.03
R4489 avss.t69 avss.n39 1271.1
R4490 avss.n806 avss.n805 1271.01
R4491 avss.n1140 avss.n87 1254.4
R4492 avss.n815 avss.n814 1251.29
R4493 avss.n520 avss.n512 1216.76
R4494 avss.n532 avss.n520 1216.76
R4495 avss.n532 avss.n531 1216.76
R4496 avss.n521 avss.n513 1216.76
R4497 avss.n524 avss.n521 1216.76
R4498 avss.n524 avss.n195 1216.76
R4499 avss.n739 avss.n734 1216.76
R4500 avss.n743 avss.n735 1216.76
R4501 avss.n903 avss.n902 1198.69
R4502 avss.n902 avss.n899 1198.69
R4503 avss.n910 avss.n905 1198.69
R4504 avss.n910 avss.n900 1198.69
R4505 avss.n1075 avss.n1074 1172.15
R4506 avss.n919 avss.n894 1167.05
R4507 avss.n901 avss.n894 1167.05
R4508 avss.n543 avss.n542 1141.23
R4509 avss.n606 avss.n603 1132.83
R4510 avss.n625 avss.n603 1132.83
R4511 avss.n612 avss.n611 1132.83
R4512 avss.n611 avss.n236 1132.83
R4513 avss.n542 avss.n541 1120.97
R4514 avss.n882 avss.n223 1100.88
R4515 avss.n883 avss.n882 1100.88
R4516 avss.n201 avss.n196 1100.88
R4517 avss.n931 avss.n196 1100.88
R4518 avss.n531 avss.n526 1100.88
R4519 avss.n526 avss.n195 1100.88
R4520 avss.n535 avss.n520 1100.88
R4521 avss.n535 avss.n521 1100.88
R4522 avss.n210 avss.n192 1100.88
R4523 avss.n210 avss.n189 1100.88
R4524 avss.n763 avss.n756 1100.88
R4525 avss.n763 avss.n751 1100.88
R4526 avss.n755 avss.n750 1100.88
R4527 avss.n791 avss.n750 1100.88
R4528 avss.n796 avss.n740 1100.88
R4529 avss.n796 avss.n746 1100.88
R4530 avss.n742 avss.n739 1100.88
R4531 avss.n743 avss.n742 1100.88
R4532 avss.n781 avss.n766 1100.88
R4533 avss.n781 avss.n769 1100.88
R4534 avss.n1083 avss.n1079 1075.2
R4535 avss.n1041 avss.n1031 1045.38
R4536 avss.n173 avss.n160 1033.74
R4537 avss.n1192 avss.n40 1032.48
R4538 avss.t19 avss.t20 1000.19
R4539 avss.t69 avss.t20 1000.19
R4540 avss.n1082 avss.n1081 999.399
R4541 avss.n626 avss.n625 994.518
R4542 avss.n626 avss.n236 994.518
R4543 avss.n628 avss.n236 994.518
R4544 avss.n616 avss.n606 994.518
R4545 avss.n616 avss.n612 994.518
R4546 avss.n614 avss.n612 994.518
R4547 avss.n573 avss.n554 994.518
R4548 avss.n574 avss.n573 994.518
R4549 avss.n574 avss.n566 994.518
R4550 avss.n566 avss.n563 994.518
R4551 avss.n592 avss.n557 994.518
R4552 avss.n567 avss.n557 994.518
R4553 avss.n568 avss.n567 994.518
R4554 avss.n568 avss.n564 994.518
R4555 avss.n621 avss.n620 981.826
R4556 dvss avss.n732 977.779
R4557 avss.n1088 avss.n1087 963.431
R4558 avss.n1085 avss.n1084 926.37
R4559 avss.n890 avss.n220 922.37
R4560 avss.n223 avss.n221 915.471
R4561 avss.n888 avss.n223 915.471
R4562 avss.n883 avss.n880 915.471
R4563 avss.n884 avss.n883 915.471
R4564 avss.n531 avss.n530 915.471
R4565 avss.n530 avss.n201 915.471
R4566 avss.n932 avss.n195 915.471
R4567 avss.n932 avss.n931 915.471
R4568 avss.n799 avss.n739 915.471
R4569 avss.n799 avss.n740 915.471
R4570 avss.n758 avss.n740 915.471
R4571 avss.n758 avss.n755 915.471
R4572 avss.n788 avss.n755 915.471
R4573 avss.n788 avss.n756 915.471
R4574 avss.n744 avss.n743 915.471
R4575 avss.n746 avss.n744 915.471
R4576 avss.n792 avss.n746 915.471
R4577 avss.n792 avss.n791 915.471
R4578 avss.n791 avss.n790 915.471
R4579 avss.n790 avss.n751 915.471
R4580 avss.t49 avss.n39 912.745
R4581 avss.t49 avss.n1175 912.745
R4582 avss.t48 avss.n1175 912.745
R4583 avss.t48 avss.n1176 912.745
R4584 avss.t18 avss.n1176 912.745
R4585 avss.t18 avss.n1192 912.745
R4586 avss.n171 avss.n169 901.063
R4587 avss.n1120 avss.n1119 882.553
R4588 avss.n1121 avss.n1120 882.553
R4589 avss.n1118 avss.n98 882.553
R4590 avss.n1122 avss.n98 882.553
R4591 avss.n623 avss.n602 881.095
R4592 avss.n1179 avss.n1177 869.38
R4593 avss.n1179 avss.n1173 869.38
R4594 avss.n1188 avss.n1178 869.38
R4595 avss.n1188 avss.n1174 869.38
R4596 avss.n1101 avss.n127 869.38
R4597 avss.n1101 avss.n128 869.38
R4598 avss.n579 avss.n566 869.38
R4599 avss.n579 avss.n568 869.38
R4600 avss.n573 avss.n572 869.38
R4601 avss.n572 avss.n557 869.38
R4602 avss.n921 avss.n920 857.888
R4603 avss.n920 avss.n919 853.793
R4604 avss.n135 avss.t66 834.323
R4605 avss.n913 avss.n899 833.155
R4606 avss.n913 avss.n900 833.155
R4607 avss.n904 avss.n903 833.155
R4608 avss.n905 avss.n904 833.155
R4609 avss.n812 avss.n811 830.769
R4610 avss.n1100 avss.t66 829.418
R4611 avss.n1100 avss.t36 829.418
R4612 avss.n1035 avss.n1032 818.081
R4613 avss.n1184 avss.n1173 734.362
R4614 avss.n1200 avss.n1173 734.362
R4615 avss.n1200 avss.n1174 734.362
R4616 avss.n1194 avss.n1174 734.362
R4617 avss.n1185 avss.n1177 734.362
R4618 avss.n1199 avss.n1177 734.362
R4619 avss.n1199 avss.n1178 734.362
R4620 avss.n1195 avss.n1178 734.362
R4621 avss.n129 avss.n127 734.362
R4622 avss.n1099 avss.n127 734.362
R4623 avss.n130 avss.n128 734.362
R4624 avss.n1094 avss.n128 734.362
R4625 avss.n658 dvss 719.574
R4626 avss.n1137 avss.n92 717.898
R4627 avss.n1130 avss.n92 717.898
R4628 avss.n1136 avss.n95 717.898
R4629 avss.n1132 avss.n95 717.898
R4630 avss.n625 avss.n624 701.432
R4631 avss.n620 avss.n606 701.432
R4632 avss.n397 avss.n268 692.46
R4633 avss.n391 avss.n268 692.46
R4634 avss.n391 avss.n390 692.46
R4635 avss.n390 avss.n389 692.46
R4636 avss.n389 avss.n274 692.46
R4637 avss.n383 avss.n274 692.46
R4638 avss.n383 avss.n382 692.46
R4639 avss.n382 avss.n381 692.46
R4640 avss.n381 avss.n281 692.46
R4641 avss.n375 avss.n281 692.46
R4642 avss.n375 avss.n374 692.46
R4643 avss.n374 avss.n373 692.46
R4644 avss.n373 avss.n293 692.46
R4645 avss.n367 avss.n293 692.46
R4646 avss.n367 avss.n366 692.46
R4647 avss.n366 avss.n365 692.46
R4648 avss.n365 avss.n305 692.46
R4649 avss.n359 avss.n305 692.46
R4650 avss.n359 avss.n358 692.46
R4651 avss.n358 avss.n357 692.46
R4652 avss.n357 avss.n317 692.46
R4653 avss.n351 avss.n317 692.46
R4654 avss.n351 avss.n350 692.46
R4655 avss.n350 avss.n349 692.46
R4656 avss.n349 avss.n329 692.46
R4657 avss.n343 avss.n329 692.46
R4658 avss.n343 avss.n342 692.46
R4659 avss.n889 avss.n222 674.668
R4660 avss.n222 avss.n216 674.668
R4661 avss.n810 avss.n809 652.436
R4662 avss.n815 avss.n810 652.436
R4663 avss.n1073 avss.n1072 640.631
R4664 avss.n171 avss.n168 639.551
R4665 avss.n593 avss.n555 636.703
R4666 avss.n565 avss.n555 636.703
R4667 avss.n580 avss.n565 636.703
R4668 avss.n581 avss.n580 636.703
R4669 avss.t9 avss.n111 634.548
R4670 avss.t1 avss.n101 634.548
R4671 avss.n583 avss.n500 632.487
R4672 avss.t9 avss.n100 622.928
R4673 avss.t1 avss.n100 622.928
R4674 avss.n627 avss.n602 622.496
R4675 avss.n1144 avss.n87 620.308
R4676 avss.t19 avss.n72 619.458
R4677 avss.n1089 avss.n158 616.385
R4678 avss.n677 avss.n218 611.778
R4679 avss.n732 avss.n731 611.778
R4680 avss.n873 avss.n219 611.778
R4681 avss.n813 avss.n652 611.778
R4682 avss.n545 avss.n510 594.447
R4683 avss.n600 avss.n599 594.447
R4684 avss.n400 avss.n399 591.17
R4685 avss.n396 avss.n395 591.169
R4686 avss.n397 avss.n396 585
R4687 avss.n270 avss.n269 585
R4688 avss.n269 avss.n268 585
R4689 avss.n393 avss.n392 585
R4690 avss.n392 avss.n391 585
R4691 avss.n273 avss.n272 585
R4692 avss.n390 avss.n273 585
R4693 avss.n388 avss.n387 585
R4694 avss.n389 avss.n388 585
R4695 avss.n386 avss.n275 585
R4696 avss.n275 avss.n274 585
R4697 avss.n385 avss.n384 585
R4698 avss.n384 avss.n383 585
R4699 avss.n280 avss.n279 585
R4700 avss.n382 avss.n280 585
R4701 avss.n380 avss.n379 585
R4702 avss.n381 avss.n380 585
R4703 avss.n378 avss.n282 585
R4704 avss.n282 avss.n281 585
R4705 avss.n377 avss.n376 585
R4706 avss.n376 avss.n375 585
R4707 avss.n292 avss.n291 585
R4708 avss.n374 avss.n292 585
R4709 avss.n372 avss.n371 585
R4710 avss.n373 avss.n372 585
R4711 avss.n370 avss.n294 585
R4712 avss.n294 avss.n293 585
R4713 avss.n369 avss.n368 585
R4714 avss.n368 avss.n367 585
R4715 avss.n304 avss.n303 585
R4716 avss.n366 avss.n304 585
R4717 avss.n364 avss.n363 585
R4718 avss.n365 avss.n364 585
R4719 avss.n362 avss.n306 585
R4720 avss.n306 avss.n305 585
R4721 avss.n361 avss.n360 585
R4722 avss.n360 avss.n359 585
R4723 avss.n316 avss.n315 585
R4724 avss.n358 avss.n316 585
R4725 avss.n356 avss.n355 585
R4726 avss.n357 avss.n356 585
R4727 avss.n354 avss.n318 585
R4728 avss.n318 avss.n317 585
R4729 avss.n353 avss.n352 585
R4730 avss.n352 avss.n351 585
R4731 avss.n328 avss.n327 585
R4732 avss.n350 avss.n328 585
R4733 avss.n348 avss.n347 585
R4734 avss.n349 avss.n348 585
R4735 avss.n346 avss.n330 585
R4736 avss.n330 avss.n329 585
R4737 avss.n345 avss.n344 585
R4738 avss.n344 avss.n343 585
R4739 avss.n341 avss.n340 585
R4740 avss.n342 avss.n341 585
R4741 avss.n399 avss.n398 585
R4742 avss.n402 avss.n401 585
R4743 avss.n403 avss.n402 585
R4744 avss.n267 avss.n266 585
R4745 avss.n404 avss.n267 585
R4746 avss.n408 avss.n407 585
R4747 avss.n407 avss.n406 585
R4748 avss.n264 avss.n263 585
R4749 avss.n405 avss.n263 585
R4750 avss.n414 avss.n413 585
R4751 avss.n414 avss.n262 585
R4752 avss.n415 avss.n260 585
R4753 avss.n416 avss.n415 585
R4754 avss.n421 avss.n261 585
R4755 avss.n417 avss.n261 585
R4756 avss.n420 avss.n419 585
R4757 avss.n419 avss.n418 585
R4758 avss.n257 avss.n256 585
R4759 avss.n256 avss.n255 585
R4760 avss.n433 avss.n432 585
R4761 avss.n434 avss.n433 585
R4762 avss.n254 avss.n253 585
R4763 avss.n435 avss.n254 585
R4764 avss.n438 avss.n437 585
R4765 avss.n437 avss.n436 585
R4766 avss.n250 avss.n249 585
R4767 avss.n249 avss.n248 585
R4768 avss.n446 avss.n445 585
R4769 avss.n447 avss.n446 585
R4770 avss.n247 avss.n246 585
R4771 avss.n448 avss.n247 585
R4772 avss.n451 avss.n450 585
R4773 avss.n450 avss.n449 585
R4774 avss.n243 avss.n241 585
R4775 avss.n241 avss.n239 585
R4776 avss.n497 avss.n496 585
R4777 avss.n498 avss.n497 585
R4778 avss.n244 avss.n242 585
R4779 avss.n242 avss.n240 585
R4780 avss.n468 avss.n467 585
R4781 avss.n468 avss.n466 585
R4782 avss.n469 avss.n458 585
R4783 avss.n470 avss.n469 585
R4784 avss.n489 avss.n459 585
R4785 avss.n471 avss.n459 585
R4786 avss.n488 avss.n460 585
R4787 avss.n472 avss.n460 585
R4788 avss.n473 avss.n461 585
R4789 avss.n474 avss.n473 585
R4790 avss.n482 avss.n464 585
R4791 avss.n475 avss.n464 585
R4792 avss.n481 avss.n465 585
R4793 avss.n476 avss.n465 585
R4794 avss.n480 avss.n478 585
R4795 avss.n478 avss.n477 585
R4796 avss.n1212 avss.t3 580.571
R4797 avss.n1222 avss.n1221 576
R4798 avss.t3 avss.n55 569.938
R4799 avss.n1218 avss.t7 559.304
R4800 avss.t7 avss.n1217 559.304
R4801 avss.n510 avss.n509 554.4
R4802 avss.n599 avss.n598 554.201
R4803 avss.n594 avss.n553 543.939
R4804 avss.n396 avss.n269 539.294
R4805 avss.n392 avss.n269 539.294
R4806 avss.n392 avss.n273 539.294
R4807 avss.n388 avss.n273 539.294
R4808 avss.n388 avss.n275 539.294
R4809 avss.n384 avss.n275 539.294
R4810 avss.n384 avss.n280 539.294
R4811 avss.n380 avss.n280 539.294
R4812 avss.n380 avss.n282 539.294
R4813 avss.n376 avss.n282 539.294
R4814 avss.n376 avss.n292 539.294
R4815 avss.n372 avss.n292 539.294
R4816 avss.n372 avss.n294 539.294
R4817 avss.n368 avss.n294 539.294
R4818 avss.n368 avss.n304 539.294
R4819 avss.n364 avss.n304 539.294
R4820 avss.n364 avss.n306 539.294
R4821 avss.n360 avss.n306 539.294
R4822 avss.n360 avss.n316 539.294
R4823 avss.n356 avss.n316 539.294
R4824 avss.n356 avss.n318 539.294
R4825 avss.n352 avss.n318 539.294
R4826 avss.n352 avss.n328 539.294
R4827 avss.n348 avss.n328 539.294
R4828 avss.n348 avss.n330 539.294
R4829 avss.n344 avss.n330 539.294
R4830 avss.n344 avss.n341 539.294
R4831 avss.n402 avss.n399 539.294
R4832 avss.n402 avss.n267 539.294
R4833 avss.n407 avss.n267 539.294
R4834 avss.n407 avss.n263 539.294
R4835 avss.n414 avss.n263 539.294
R4836 avss.n415 avss.n414 539.294
R4837 avss.n415 avss.n261 539.294
R4838 avss.n419 avss.n261 539.294
R4839 avss.n419 avss.n256 539.294
R4840 avss.n433 avss.n256 539.294
R4841 avss.n433 avss.n254 539.294
R4842 avss.n437 avss.n254 539.294
R4843 avss.n437 avss.n249 539.294
R4844 avss.n446 avss.n249 539.294
R4845 avss.n446 avss.n247 539.294
R4846 avss.n450 avss.n247 539.294
R4847 avss.n450 avss.n241 539.294
R4848 avss.n497 avss.n241 539.294
R4849 avss.n497 avss.n242 539.294
R4850 avss.n468 avss.n242 539.294
R4851 avss.n469 avss.n468 539.294
R4852 avss.n469 avss.n459 539.294
R4853 avss.n460 avss.n459 539.294
R4854 avss.n473 avss.n460 539.294
R4855 avss.n473 avss.n464 539.294
R4856 avss.n465 avss.n464 539.294
R4857 avss.n478 avss.n465 539.294
R4858 avss.n1064 avss.n176 538.484
R4859 avss.n1070 avss.n176 538.484
R4860 avss.n24 avss.n10 538.038
R4861 avss.n922 avss.n200 535.072
R4862 avss.n1208 avss.n1206 532.726
R4863 avss.n912 avss.n901 518.009
R4864 avss.n912 avss.n911 518.009
R4865 avss.n783 avss.n754 515.035
R4866 avss.n783 avss.n782 515.035
R4867 avss.n782 avss.n768 515.035
R4868 avss.n814 avss.n175 510.603
R4869 avss.t63 avss.n116 506.709
R4870 avss.n1061 avss.n183 479.248
R4871 avss.n602 avss.n500 476.474
R4872 avss.n101 avss.n93 474.168
R4873 avss.n805 avss.n733 466.197
R4874 avss.n741 avss.n733 466.197
R4875 avss.t32 avss.n9 463.606
R4876 avss.t32 avss.n10 463.606
R4877 avss.t52 avss.n94 463.606
R4878 avss.n94 avss.t53 463.606
R4879 avss.t52 avss.n93 454.515
R4880 avss.n118 avss.n117 443.952
R4881 avss.n1085 avss.n163 443.057
R4882 avss.n1213 avss.n1212 442.339
R4883 avss.n1222 avss.n50 440.32
R4884 avss.n541 avss.n511 429.568
R4885 avss.n534 avss.n511 429.568
R4886 avss.n534 avss.n533 429.568
R4887 avss.n1037 avss.n1036 426.846
R4888 avss.n117 avss.n111 402.113
R4889 avss.n1209 avss.n1208 401.372
R4890 avss.n470 avss.n466 390.029
R4891 avss.n471 avss.n470 390.029
R4892 avss.n472 avss.n471 390.029
R4893 avss.n474 avss.n472 390.029
R4894 avss.n475 avss.n474 390.029
R4895 avss.n476 avss.n475 390.029
R4896 avss.n477 avss.n476 390.029
R4897 avss.n1257 avss.n6 387.457
R4898 avss.n1206 avss.n62 381.137
R4899 avss.t65 avss.n72 380.731
R4900 avss.n466 avss.n240 379.801
R4901 avss.n403 avss.n398 371.505
R4902 avss.n404 avss.n403 371.505
R4903 avss.n406 avss.n404 371.505
R4904 avss.n406 avss.n405 371.505
R4905 avss.n405 avss.n262 371.505
R4906 avss.n416 avss.n262 371.505
R4907 avss.n417 avss.n416 371.505
R4908 avss.n418 avss.n417 371.505
R4909 avss.n418 avss.n255 371.505
R4910 avss.n434 avss.n255 371.505
R4911 avss.n435 avss.n434 371.505
R4912 avss.n436 avss.n435 371.505
R4913 avss.n436 avss.n248 371.505
R4914 avss.n447 avss.n248 371.505
R4915 avss.n448 avss.n447 371.505
R4916 avss.n449 avss.n448 371.505
R4917 avss.n449 avss.n239 371.505
R4918 avss.n498 avss.n240 371.505
R4919 avss.n1096 avss.n1091 370.957
R4920 avss.t5 avss.n24 367.908
R4921 avss.t5 avss.n1256 367.908
R4922 avss.n602 avss.n217 363.445
R4923 avss.n582 avss.n581 360.517
R4924 avss.n917 avss.n897 356.142
R4925 avss.n798 avss.n741 350.757
R4926 avss.n798 avss.n797 350.757
R4927 avss.n797 avss.n745 350.757
R4928 avss.n753 avss.n745 350.757
R4929 avss.n789 avss.n753 350.757
R4930 avss.n789 avss.n754 350.757
R4931 avss.n173 avss.n136 348.188
R4932 avss.n908 avss.n183 337.695
R4933 avss.n213 avss.n212 335.473
R4934 avss.n1217 avss.n9 325.375
R4935 avss.n814 avss.n813 324.808
R4936 avss.n1087 avss.n160 321.82
R4937 avss.n211 avss.n191 315.017
R4938 avss.t13 avss.n40 314.741
R4939 avss.t0 avss.n1213 314.741
R4940 avss.n1209 avss.n5 313.601
R4941 avss.n525 avss.n190 310.925
R4942 avss.n1110 avss.n110 304.849
R4943 avss.n150 avss.n149 302.017
R4944 dvss avss.n659 301.029
R4945 avss.n499 avss.n498 297.978
R4946 avss.n78 avss.n64 292.5
R4947 avss.n78 avss.t59 292.5
R4948 avss.n75 avss.n31 292.5
R4949 avss.t59 avss.n75 292.5
R4950 avss.n790 avss.n752 292.5
R4951 avss.n790 avss.n789 292.5
R4952 avss.n793 avss.n792 292.5
R4953 avss.n792 avss.n745 292.5
R4954 avss.n748 avss.n744 292.5
R4955 avss.n798 avss.n744 292.5
R4956 avss.n800 avss.n799 292.5
R4957 avss.n799 avss.n798 292.5
R4958 avss.n759 avss.n758 292.5
R4959 avss.n758 avss.n745 292.5
R4960 avss.n788 avss.n787 292.5
R4961 avss.n789 avss.n788 292.5
R4962 avss.n817 avss.n816 292.5
R4963 avss.n816 avss.n815 292.5
R4964 avss.n808 avss.n807 292.5
R4965 avss.n809 avss.n808 292.5
R4966 avss.n933 avss.n932 292.5
R4967 avss.n932 avss.n191 292.5
R4968 avss.n530 avss.n529 292.5
R4969 avss.n530 avss.n191 292.5
R4970 avss.n885 avss.n884 292.5
R4971 avss.n884 avss.n216 292.5
R4972 avss.n880 avss.n879 292.5
R4973 avss.n880 avss.n216 292.5
R4974 avss.n228 avss.n221 292.5
R4975 avss.n889 avss.n221 292.5
R4976 avss.n888 avss.n887 292.5
R4977 avss.n889 avss.n888 292.5
R4978 avss.n726 avss.n723 292.443
R4979 avss.n158 avss.t15 291.185
R4980 avss.n1064 avss.n1063 286.646
R4981 avss.n583 avss.n582 276.187
R4982 avss.n1246 avss.n27 274.389
R4983 avss.n150 avss.t15 266.839
R4984 avss.n1095 avss.n116 262.652
R4985 avss.n549 avss.n548 252.941
R4986 avss.n596 avss.n504 252.941
R4987 avss.n613 avss.n235 247.719
R4988 avss.n1146 avss.n80 244.329
R4989 avss.n1151 avss.n80 244.329
R4990 avss.n1155 avss.n1154 244.329
R4991 avss.n1154 avss.n1153 244.329
R4992 avss.n1239 avss.n35 244.329
R4993 avss.n1239 avss.n1238 244.329
R4994 avss.n892 avss.n217 241.185
R4995 avss.n1139 avss.n89 227.097
R4996 avss.n1128 avss.n1126 216.847
R4997 avss.n906 avss.n897 214.589
R4998 avss.n619 avss.n607 214.213
R4999 avss.n1253 avss.n1252 211.93
R5000 avss.n1061 avss.n1060 210.745
R5001 avss.n1134 avss.n1126 210.447
R5002 avss.n1218 avss.n1215 206.284
R5003 avss.n1068 avss.n179 202.918
R5004 avss.n1068 avss.n1067 202.918
R5005 avss.n1067 avss.n1066 202.918
R5006 avss.n1066 avss.n179 202.918
R5007 avss.t5 avss.n1257 195
R5008 avss.n1259 avss.n1258 195
R5009 avss.n1258 avss.t5 195
R5010 avss.t47 avss.t44 191.756
R5011 avss.t12 avss.t47 191.756
R5012 avss.t30 avss.t12 191.756
R5013 avss.t61 avss.t30 191.756
R5014 avss.t74 avss.t61 191.756
R5015 avss.t41 avss.t74 191.756
R5016 avss.t41 avss.t28 191.756
R5017 avss.t28 avss.t71 191.756
R5018 avss.t44 avss.t46 191.526
R5019 avss.n1186 avss.n1181 187.859
R5020 avss.n1196 avss.n1190 187.859
R5021 avss.n1265 avss.n5 186.058
R5022 avss.n917 avss.n916 181.679
R5023 avss.n813 dvss 181.288
R5024 avss.n1111 avss.n119 177.589
R5025 avss.t70 avss.t39 175.409
R5026 avss.t39 avss.t58 175.409
R5027 avss.t58 avss.t72 175.409
R5028 avss.t25 avss.n41 170.815
R5029 avss.t35 avss.n41 170.815
R5030 avss.n149 avss.t46 170.606
R5031 avss.t71 avss.t68 165.79
R5032 avss.n1183 avss.n1181 165.014
R5033 avss.n1193 avss.n1190 165.014
R5034 avss.n1242 avss.t20 164.179
R5035 avss.n936 avss.n190 163.645
R5036 avss.n142 avss.n30 161.438
R5037 avss.n936 avss.n191 159.554
R5038 avss.n778 avss.n772 159.054
R5039 avss.n927 avss.n926 159.011
R5040 avss.n1255 avss.t72 156.388
R5041 avss.n803 avss.n736 150.399
R5042 avss.n539 avss.n538 150.398
R5043 avss.t68 avss.t60 147.317
R5044 avss.t16 avss.t29 147.317
R5045 avss.t75 avss.t38 147.317
R5046 avss.t43 avss.t62 147.317
R5047 avss.t62 avss.t40 147.317
R5048 avss.t40 avss.t26 147.317
R5049 avss.t26 avss.t42 147.317
R5050 avss.t42 avss.t54 147.317
R5051 avss.t54 avss.t22 147.317
R5052 avss.t22 avss.t34 147.317
R5053 avss.t34 avss.t51 147.317
R5054 avss.t51 avss.t55 147.317
R5055 avss.t55 avss.t21 147.317
R5056 avss.t23 avss.t56 147.317
R5057 avss.n1262 avss.n1261 146.25
R5058 avss.t32 avss.n1262 146.25
R5059 avss.n1264 avss.n1263 146.25
R5060 avss.n1263 avss.t32 146.25
R5061 avss.n1196 avss.n1195 146.25
R5062 avss.n1195 avss.t18 146.25
R5063 avss.n1199 avss.n1198 146.25
R5064 avss.t48 avss.n1199 146.25
R5065 avss.n1186 avss.n1185 146.25
R5066 avss.n1185 avss.t49 146.25
R5067 avss.n1194 avss.n1193 146.25
R5068 avss.t18 avss.n1194 146.25
R5069 avss.n1201 avss.n1200 146.25
R5070 avss.n1200 avss.t48 146.25
R5071 avss.n1184 avss.n1183 146.25
R5072 avss.t49 avss.n1184 146.25
R5073 avss.n776 avss.n772 146.25
R5074 avss.n776 avss.n775 146.25
R5075 avss.n742 avss.n737 146.25
R5076 avss.n742 avss.n741 146.25
R5077 avss.n796 avss.n795 146.25
R5078 avss.n797 avss.n796 146.25
R5079 avss.n757 avss.n750 146.25
R5080 avss.n753 avss.n750 146.25
R5081 avss.n764 avss.n763 146.25
R5082 avss.n763 avss.n754 146.25
R5083 avss.n781 avss.n780 146.25
R5084 avss.n782 avss.n781 146.25
R5085 avss.n736 avss.n735 146.25
R5086 avss.n735 avss.n733 146.25
R5087 avss.n804 avss.n803 146.25
R5088 avss.n805 avss.n804 146.25
R5089 avss.n802 avss.n734 146.25
R5090 avss.n734 avss.n733 146.25
R5091 avss.n657 avss.n655 146.25
R5092 avss.n810 avss.n657 146.25
R5093 avss.n656 avss.n654 146.25
R5094 avss.n810 avss.n656 146.25
R5095 avss.n545 avss.n544 146.25
R5096 avss.n544 avss.n543 146.25
R5097 avss.n550 avss.n549 146.25
R5098 avss.n551 avss.n550 146.25
R5099 avss.n596 avss.n595 146.25
R5100 avss.n595 avss.n594 146.25
R5101 avss.n601 avss.n600 146.25
R5102 avss.n620 avss.n619 146.25
R5103 avss.n624 avss.n605 146.25
R5104 avss.n624 avss.n623 146.25
R5105 avss.n210 avss.n209 146.25
R5106 avss.n211 avss.n210 146.25
R5107 avss.n188 avss.n186 146.25
R5108 avss.n525 avss.n188 146.25
R5109 avss.n536 avss.n535 146.25
R5110 avss.n535 avss.n534 146.25
R5111 avss.n527 avss.n526 146.25
R5112 avss.n526 avss.n190 146.25
R5113 avss.n204 avss.n196 146.25
R5114 avss.n212 avss.n196 146.25
R5115 avss.n524 avss.n523 146.25
R5116 avss.n533 avss.n524 146.25
R5117 avss.n514 avss.n513 146.25
R5118 avss.n513 avss.n511 146.25
R5119 avss.n540 avss.n539 146.25
R5120 avss.n541 avss.n540 146.25
R5121 avss.n538 avss.n512 146.25
R5122 avss.n512 avss.n511 146.25
R5123 avss.n532 avss.n515 146.25
R5124 avss.n533 avss.n532 146.25
R5125 avss.n882 avss.n881 146.25
R5126 avss.n882 avss.n222 146.25
R5127 avss.n886 avss.n224 146.25
R5128 avss.n224 avss.n222 146.25
R5129 avss.n229 avss.n227 146.25
R5130 avss.n227 avss.n222 146.25
R5131 avss.n924 avss.n923 146.25
R5132 avss.n923 avss.n922 146.25
R5133 avss.n926 avss.n197 146.25
R5134 avss.n921 avss.n197 146.25
R5135 avss.n1099 avss.n1098 146.25
R5136 avss.t36 avss.n1099 146.25
R5137 avss.n131 avss.n129 146.25
R5138 avss.n129 avss.t66 146.25
R5139 avss.n1112 avss.n1111 146.25
R5140 avss.t63 avss.n1112 146.25
R5141 avss.n1138 avss.n1137 146.25
R5142 avss.n1137 avss.t52 146.25
R5143 avss.n1130 avss.n1129 146.25
R5144 avss.n1130 avss.t53 146.25
R5145 avss.n1094 avss.n1093 146.25
R5146 avss.t36 avss.n1094 146.25
R5147 avss.n132 avss.n130 146.25
R5148 avss.n130 avss.t66 146.25
R5149 avss.n1114 avss.n1113 146.25
R5150 avss.n1113 avss.t63 146.25
R5151 avss.n1133 avss.n1132 146.25
R5152 avss.n1132 avss.t53 146.25
R5153 avss.n1136 avss.n1135 146.25
R5154 avss.t52 avss.n1136 146.25
R5155 avss.n629 avss.n235 145.726
R5156 avss.t38 avss.n1231 143.768
R5157 avss.n145 avss.t45 141.994
R5158 avss.t27 avss.n85 141.994
R5159 avss.n909 avss.n908 141.554
R5160 avss.n906 avss.n898 141.554
R5161 avss.t56 avss.t70 140.431
R5162 avss.n607 avss.n605 140.059
R5163 avss.t69 avss.t31 135.781
R5164 avss.n610 avss.n234 134.024
R5165 avss.n618 avss.n609 134.024
R5166 avss.n110 avss.n109 133.369
R5167 avss.n1168 avss.n44 131.964
R5168 avss.t33 avss.n73 131.344
R5169 avss.t59 avss.n77 131.344
R5170 avss.n909 avss.n184 131.012
R5171 avss.n915 avss.n898 131.012
R5172 avss.n807 avss.n654 131.012
R5173 avss.n807 avss.n655 131.012
R5174 avss.n229 avss.n228 131.012
R5175 avss.n887 avss.n886 131.012
R5176 avss.n213 avss.n199 130.917
R5177 avss.n133 avss.n131 130.087
R5178 avss.n586 avss.n561 127.703
R5179 avss.n630 avss.n234 126.495
R5180 avss.n609 avss.n608 126.495
R5181 avss.n556 avss.n553 124.909
R5182 avss.n1215 avss.n55 123.346
R5183 avss.n1111 avss.n1110 120.472
R5184 avss.n570 avss.n569 120.088
R5185 avss.t19 avss.n1160 119.806
R5186 avss.n1237 avss.n37 119.575
R5187 avss.n1096 avss.n1095 118.919
R5188 avss.n1247 avss.n1246 118.722
R5189 avss.n533 avss.n525 118.642
R5190 avss.n58 avss.n53 117.001
R5191 avss.t7 avss.n53 117.001
R5192 avss.n54 avss.n5 117.001
R5193 avss.t7 avss.n54 117.001
R5194 avss.n57 avss.n56 117.001
R5195 avss.n56 avss.t3 117.001
R5196 avss.n1210 avss.n1209 117.001
R5197 avss.n1210 avss.t3 117.001
R5198 avss.n1237 avss.n1236 117.001
R5199 avss.n1236 avss.t69 117.001
R5200 avss.n69 avss.n36 117.001
R5201 avss.n69 avss.t20 117.001
R5202 avss.n1152 avss.n71 117.001
R5203 avss.t19 avss.n71 117.001
R5204 avss.n1150 avss.n1149 117.001
R5205 avss.n1149 avss.t65 117.001
R5206 avss.n1148 avss.n1147 117.001
R5207 avss.t65 avss.n1148 117.001
R5208 avss.n1161 avss.n68 117.001
R5209 avss.n1161 avss.t19 117.001
R5210 avss.n1164 avss.n1163 117.001
R5211 avss.n1163 avss.t20 117.001
R5212 avss.n1235 avss.n1234 117.001
R5213 avss.t69 avss.n1235 117.001
R5214 avss.n778 avss.n777 117.001
R5215 avss.n777 avss.n768 117.001
R5216 avss.n771 avss.n767 117.001
R5217 avss.n783 avss.n767 117.001
R5218 avss.n785 avss.n784 117.001
R5219 avss.n784 avss.n783 117.001
R5220 avss.n774 avss.n773 117.001
R5221 avss.n774 avss.n768 117.001
R5222 avss.n208 avss.n203 117.001
R5223 avss.n208 avss.n199 117.001
R5224 avss.n938 avss.n937 117.001
R5225 avss.n937 avss.n936 117.001
R5226 avss.n935 avss.n934 117.001
R5227 avss.n936 avss.n935 117.001
R5228 avss.n207 avss.n206 117.001
R5229 avss.n207 avss.n199 117.001
R5230 avss.n930 avss.n198 117.001
R5231 avss.n930 avss.n929 117.001
R5232 avss.n928 avss.n927 117.001
R5233 avss.n929 avss.n928 117.001
R5234 avss.n907 avss.n904 117.001
R5235 avss.n912 avss.n904 117.001
R5236 avss.n914 avss.n913 117.001
R5237 avss.n913 avss.n912 117.001
R5238 avss.n179 avss.n177 117.001
R5239 avss.n177 avss.n176 117.001
R5240 avss.n1067 avss.n178 117.001
R5241 avss.n178 avss.n176 117.001
R5242 avss.n139 avss.n137 117.001
R5243 avss.n137 avss.t15 117.001
R5244 avss.n155 avss.n138 117.001
R5245 avss.n138 avss.t15 117.001
R5246 avss.n1121 avss.n89 117.001
R5247 avss.t1 avss.n1121 117.001
R5248 avss.n1119 avss.n110 117.001
R5249 avss.n1119 avss.t9 117.001
R5250 avss.n1123 avss.n1122 117.001
R5251 avss.n1122 avss.t1 117.001
R5252 avss.n1118 avss.n1117 117.001
R5253 avss.t9 avss.n1118 117.001
R5254 avss.n618 avss.n617 113.695
R5255 avss.n617 avss.n610 113.695
R5256 avss.n613 avss.n610 113.695
R5257 avss.n571 avss.n570 113.695
R5258 avss.n575 avss.n571 113.695
R5259 avss.n576 avss.n575 113.695
R5260 avss.n576 avss.n561 113.695
R5261 avss.n924 avss.n203 110.438
R5262 avss.n1233 avss.n28 108.906
R5263 avss.n732 dvss 108.642
R5264 avss.n1098 avss.n125 105.412
R5265 avss.n1197 avss.n1189 103.906
R5266 avss.n1187 avss.n1180 103.906
R5267 avss.n571 avss.n559 103.906
R5268 avss.n578 avss.n576 103.906
R5269 avss.n1265 avss.n1264 103.772
R5270 avss.n1264 avss.n6 101.944
R5271 avss.n590 avss.n559 101.647
R5272 avss.n578 avss.n577 101.647
R5273 avss.n1189 avss.n1172 100.141
R5274 avss.n1180 avss.n1171 100.141
R5275 avss.t21 avss.t13 99.3954
R5276 avss.n929 avss.n200 98.1874
R5277 avss.n1182 avss.n1181 97.5005
R5278 avss.n1182 avss.n39 97.5005
R5279 avss.n1180 avss.n1179 97.5005
R5280 avss.n1179 avss.n1175 97.5005
R5281 avss.n1189 avss.n1188 97.5005
R5282 avss.n1188 avss.n1176 97.5005
R5283 avss.n1191 avss.n1190 97.5005
R5284 avss.n1192 avss.n1191 97.5005
R5285 avss.n585 avss.n584 97.5005
R5286 avss.n584 avss.n583 97.5005
R5287 avss.n572 avss.n559 97.5005
R5288 avss.n572 avss.n555 97.5005
R5289 avss.n563 avss.n561 97.5005
R5290 avss.n581 avss.n563 97.5005
R5291 avss.n575 avss.n574 97.5005
R5292 avss.n574 avss.n565 97.5005
R5293 avss.n570 avss.n554 97.5005
R5294 avss.n593 avss.n554 97.5005
R5295 avss.n579 avss.n578 97.5005
R5296 avss.n580 avss.n579 97.5005
R5297 avss.n564 avss.n562 97.5005
R5298 avss.n581 avss.n564 97.5005
R5299 avss.n567 avss.n560 97.5005
R5300 avss.n567 avss.n565 97.5005
R5301 avss.n592 avss.n591 97.5005
R5302 avss.n593 avss.n592 97.5005
R5303 avss.n569 avss.n556 97.5005
R5304 avss.n614 avss.n613 97.5005
R5305 avss.n615 avss.n614 97.5005
R5306 avss.n617 avss.n616 97.5005
R5307 avss.n616 avss.n615 97.5005
R5308 avss.n629 avss.n628 97.5005
R5309 avss.n628 avss.n627 97.5005
R5310 avss.n626 avss.n233 97.5005
R5311 avss.n627 avss.n626 97.5005
R5312 avss.n1066 avss.n1065 97.5005
R5313 avss.n1065 avss.n1064 97.5005
R5314 avss.n1069 avss.n1068 97.5005
R5315 avss.n1070 avss.n1069 97.5005
R5316 avss.n134 avss.n133 97.5005
R5317 avss.n135 avss.n134 97.5005
R5318 avss.n1102 avss.n1101 97.5005
R5319 avss.n1101 avss.n1100 97.5005
R5320 avss.n1097 avss.n124 97.5005
R5321 avss.n1097 avss.n1096 97.5005
R5322 avss.n59 avss.n57 97.4474
R5323 avss.n57 avss.n45 96.377
R5324 avss.n1160 avss.n74 95.8456
R5325 avss.n907 avss.n906 95.2476
R5326 avss.n908 avss.n907 95.2476
R5327 avss.n142 avss.n141 92.9825
R5328 avss.n773 avss.n772 92.4525
R5329 avss.n939 avss.n186 91.8104
R5330 avss.n817 avss.n655 90.905
R5331 avss.n1232 avss.t75 90.5209
R5332 avss.n803 avss.n802 90.4228
R5333 avss.n1143 avss.n1142 89.1641
R5334 avss.n1233 avss.n37 88.375
R5335 avss.n1115 avss.n112 87.9969
R5336 avss.n109 avss.n89 87.9489
R5337 avss.n818 avss.n654 87.6306
R5338 avss.n771 avss.n770 87.3417
R5339 avss.n779 avss.n771 87.3417
R5340 avss.n779 avss.n778 87.3417
R5341 avss.n927 avss.n202 87.3417
R5342 avss.n539 avss.n514 86.4517
R5343 avss.n1098 avss.n124 85.4292
R5344 avss.n119 avss.n113 84.8377
R5345 avss.n1187 avss.n1186 83.9534
R5346 avss.n1198 avss.n1187 83.9534
R5347 avss.n1198 avss.n1197 83.9534
R5348 avss.n1197 avss.n1196 83.9534
R5349 avss.n1079 avss.n1078 83.7224
R5350 avss.n1141 avss.n1140 83.407
R5351 avss.n1170 avss.t50 83.0379
R5352 avss.n1145 avss.n1144 81.6649
R5353 avss.n1261 avss.n1260 81.2016
R5354 avss.n1127 avss.n81 80.6409
R5355 avss.n619 avss.n618 80.1887
R5356 avss.n1241 avss.t31 79.8714
R5357 avss.n879 avss.n229 79.57
R5358 avss.n886 avss.n885 79.57
R5359 avss.n747 avss.n736 79.0593
R5360 avss.n538 avss.n537 79.0593
R5361 avss.n537 avss.n515 79.0593
R5362 avss.n528 avss.n515 79.0593
R5363 avss.t19 avss.n73 78.984
R5364 avss.n124 avss.t37 78.1972
R5365 avss.n1102 avss.t67 78.1972
R5366 avss.n1060 avss.n1059 75.8227
R5367 avss.n156 avss.n139 75.4543
R5368 avss.t65 avss.t45 73.6592
R5369 avss.t65 avss.t27 73.6592
R5370 avss.n1229 avss.t25 73.6592
R5371 avss.n499 avss.n239 73.5273
R5372 avss.n926 avss.n925 73.0738
R5373 avss.n925 avss.n924 72.206
R5374 avss.n204 avss.n202 71.5299
R5375 avss.n205 avss.n204 71.5299
R5376 avss.n786 avss.n764 71.5299
R5377 avss.n770 avss.n764 71.5299
R5378 avss.n760 avss.n757 71.5299
R5379 avss.n757 avss.n749 71.5299
R5380 avss.n795 avss.n738 71.5299
R5381 avss.n795 avss.n794 71.5299
R5382 avss.n801 avss.n737 71.5299
R5383 avss.n747 avss.n737 71.5299
R5384 avss.n780 avss.n765 71.5299
R5385 avss.n780 avss.n779 71.5299
R5386 avss.n881 avss.n225 71.5299
R5387 avss.n209 avss.n194 71.5299
R5388 avss.n209 avss.n187 71.5299
R5389 avss.n522 avss.n186 71.5299
R5390 avss.n528 avss.n527 71.5299
R5391 avss.n527 avss.n193 71.5299
R5392 avss.n537 avss.n536 71.5299
R5393 avss.n536 avss.n519 71.5299
R5394 avss.n21 avss.n16 71.2831
R5395 avss.n881 avss.n226 70.777
R5396 avss.t65 avss.t53 70.1793
R5397 avss.n1158 avss.n1157 70.0532
R5398 avss.n1230 avss.t35 69.4486
R5399 avss.t0 avss.n1214 69.4486
R5400 avss.n141 avss.n79 69.1602
R5401 avss.n1089 avss.n1088 69.1236
R5402 avss.n1207 avss.n41 67.8493
R5403 avss.n156 avss.n155 66.6531
R5404 avss.n585 avss.n562 66.3047
R5405 avss.n65 avss.n32 65.9625
R5406 avss.n1133 avss.n1127 65.4191
R5407 avss.n594 avss.n593 65.3575
R5408 avss.n1245 avss.n1244 65.1217
R5409 avss.n1220 avss.n1219 65.0005
R5410 avss.n1219 avss.n1218 65.0005
R5411 avss.n1216 avss.n52 65.0005
R5412 avss.n1217 avss.n1216 65.0005
R5413 avss.n1208 avss.n1207 65.0005
R5414 avss.n1228 avss.n1227 65.0005
R5415 avss.n1229 avss.n1228 65.0005
R5416 avss.n607 avss.n604 65.0005
R5417 avss.n609 avss.n603 65.0005
R5418 avss.n622 avss.n603 65.0005
R5419 avss.n611 avss.n234 65.0005
R5420 avss.n611 avss.n238 65.0005
R5421 avss.n237 avss.n235 65.0005
R5422 avss.n238 avss.n237 65.0005
R5423 avss.n918 avss.n917 65.0005
R5424 avss.n919 avss.n918 65.0005
R5425 avss.n902 avss.n898 65.0005
R5426 avss.n902 avss.n901 65.0005
R5427 avss.n910 avss.n909 65.0005
R5428 avss.n911 avss.n910 65.0005
R5429 avss.n1062 avss.n1061 65.0005
R5430 avss.n1063 avss.n1062 65.0005
R5431 avss.n1183 avss.n1171 64.8732
R5432 avss.n1201 avss.n1172 64.8732
R5433 avss.n1193 avss.n1172 64.8732
R5434 avss.n1202 avss.n1171 64.2914
R5435 avss.t63 avss.n118 62.758
R5436 avss.n131 avss.n125 62.4946
R5437 avss.n1252 avss.n28 61.5624
R5438 avss.n591 avss.n558 60.3224
R5439 avss.n748 avss.n747 59.4829
R5440 avss.n794 avss.n748 59.4829
R5441 avss.n794 avss.n793 59.4829
R5442 avss.n793 avss.n749 59.4829
R5443 avss.n752 avss.n749 59.4829
R5444 avss.n770 avss.n752 59.4829
R5445 avss.n228 avss.n225 59.4829
R5446 avss.n887 avss.n225 59.4829
R5447 avss.n529 avss.n528 59.4829
R5448 avss.n529 avss.n202 59.4829
R5449 avss.n1227 avss.n1226 59.2721
R5450 avss.t29 avss.n1232 56.7976
R5451 avss.n1080 avss.n159 54.7639
R5452 avss.n1072 avss.n136 52.0595
R5453 avss.n1242 avss.n1241 51.4729
R5454 avss.n916 avss.n915 50.6672
R5455 avss.n77 avss.t20 48.8105
R5456 avss.n152 avss.n151 48.7505
R5457 avss.n151 avss.n150 48.7505
R5458 avss.n157 avss.n156 48.7505
R5459 avss.n158 avss.n157 48.7505
R5460 avss.n1226 avss.n45 48.0896
R5461 avss.t35 avss.t57 47.9231
R5462 avss.t0 avss.t23 47.9231
R5463 avss.n1131 avss.n72 46.8649
R5464 avss.n154 avss.n153 46.2264
R5465 avss.n133 avss.n132 43.5408
R5466 avss.n1249 avss.t73 42.3691
R5467 avss.n23 avss.n22 41.7862
R5468 avss.n1256 avss.n23 41.7862
R5469 avss.n49 avss.n14 41.7862
R5470 avss.n24 avss.n14 41.7862
R5471 avss.n897 avss.n895 41.7862
R5472 avss.n895 avss.n894 41.7862
R5473 avss.n916 avss.n896 41.7862
R5474 avss.n896 avss.n894 41.7862
R5475 avss.n153 avss.n86 41.5158
R5476 avss.n15 avss.n13 41.5006
R5477 avss.n1145 avss.n86 41.2882
R5478 avss.n1206 avss.t14 41.0016
R5479 avss.n1140 avss.n1139 40.465
R5480 avss.n108 avss.t2 39.0988
R5481 avss.n105 avss.t4 39.0988
R5482 avss.n1106 avss.t11 39.0988
R5483 avss.n1220 avss.t8 39.0988
R5484 avss.n120 avss.t10 39.0988
R5485 avss.n51 avss.n7 39.0005
R5486 avss.n9 avss.n7 39.0005
R5487 avss.n12 avss.n8 39.0005
R5488 avss.n10 avss.n8 39.0005
R5489 avss.n122 avss.n115 39.0005
R5490 avss.n117 avss.n115 39.0005
R5491 avss.n119 avss.n114 39.0005
R5492 avss.n116 avss.n114 39.0005
R5493 avss.n96 avss.n91 39.0005
R5494 avss.n93 avss.n91 39.0005
R5495 avss.n1126 avss.n1125 39.0005
R5496 avss.n1125 avss.n94 39.0005
R5497 avss.n1131 avss.n1127 39.0005
R5498 avss.n938 avss.n187 38.5667
R5499 avss.n203 avss.n187 38.5667
R5500 avss.n1142 avss.n87 38.4005
R5501 avss.n871 avss.n635 36.1417
R5502 avss.n866 avss.n865 36.1417
R5503 avss.n861 avss.n860 36.1417
R5504 avss.n860 avss.n859 36.1417
R5505 avss.n859 avss.n639 36.1417
R5506 avss.n855 avss.n639 36.1417
R5507 avss.n853 avss.n641 36.1417
R5508 avss.n849 avss.n641 36.1417
R5509 avss.n849 avss.n848 36.1417
R5510 avss.n848 avss.n847 36.1417
R5511 avss.n841 avss.n645 36.1417
R5512 avss.n830 avss.n829 36.1417
R5513 avss.n719 avss.n718 36.1417
R5514 avss.n713 avss.n663 36.1417
R5515 avss.n717 avss.n663 36.1417
R5516 avss.n711 avss.n665 36.1417
R5517 avss.n712 avss.n711 36.1417
R5518 avss.n699 avss.n698 36.1417
R5519 avss.n700 avss.n699 36.1417
R5520 avss.n700 avss.n668 36.1417
R5521 avss.n704 avss.n668 36.1417
R5522 avss.n688 avss.n687 36.1417
R5523 avss.n688 avss.n672 36.1417
R5524 avss.n692 avss.n672 36.1417
R5525 avss.n693 avss.n692 36.1417
R5526 avss.n694 avss.n693 36.1417
R5527 avss.n681 avss.n675 36.1417
R5528 avss.n685 avss.n675 36.1417
R5529 avss.n393 avss.n270 36.1417
R5530 avss.n393 avss.n272 36.1417
R5531 avss.n387 avss.n272 36.1417
R5532 avss.n387 avss.n386 36.1417
R5533 avss.n386 avss.n385 36.1417
R5534 avss.n385 avss.n279 36.1417
R5535 avss.n379 avss.n279 36.1417
R5536 avss.n379 avss.n378 36.1417
R5537 avss.n378 avss.n377 36.1417
R5538 avss.n377 avss.n291 36.1417
R5539 avss.n371 avss.n291 36.1417
R5540 avss.n371 avss.n370 36.1417
R5541 avss.n370 avss.n369 36.1417
R5542 avss.n369 avss.n303 36.1417
R5543 avss.n363 avss.n303 36.1417
R5544 avss.n363 avss.n362 36.1417
R5545 avss.n362 avss.n361 36.1417
R5546 avss.n361 avss.n315 36.1417
R5547 avss.n355 avss.n315 36.1417
R5548 avss.n355 avss.n354 36.1417
R5549 avss.n354 avss.n353 36.1417
R5550 avss.n353 avss.n327 36.1417
R5551 avss.n347 avss.n327 36.1417
R5552 avss.n347 avss.n346 36.1417
R5553 avss.n346 avss.n345 36.1417
R5554 avss.n345 avss.n340 36.1417
R5555 avss.n401 avss.n266 36.1417
R5556 avss.n408 avss.n266 36.1417
R5557 avss.n408 avss.n264 36.1417
R5558 avss.n413 avss.n264 36.1417
R5559 avss.n413 avss.n260 36.1417
R5560 avss.n421 avss.n260 36.1417
R5561 avss.n421 avss.n420 36.1417
R5562 avss.n420 avss.n257 36.1417
R5563 avss.n432 avss.n257 36.1417
R5564 avss.n432 avss.n253 36.1417
R5565 avss.n438 avss.n253 36.1417
R5566 avss.n438 avss.n250 36.1417
R5567 avss.n445 avss.n250 36.1417
R5568 avss.n445 avss.n246 36.1417
R5569 avss.n451 avss.n246 36.1417
R5570 avss.n451 avss.n243 36.1417
R5571 avss.n496 avss.n243 36.1417
R5572 avss.n496 avss.n244 36.1417
R5573 avss.n467 avss.n244 36.1417
R5574 avss.n467 avss.n458 36.1417
R5575 avss.n489 avss.n458 36.1417
R5576 avss.n489 avss.n488 36.1417
R5577 avss.n488 avss.n461 36.1417
R5578 avss.n482 avss.n461 36.1417
R5579 avss.n482 avss.n481 36.1417
R5580 avss.n481 avss.n480 36.1417
R5581 avss.t59 avss.n74 35.4987
R5582 avss.n698 avss.n670 35.0123
R5583 avss.n622 avss.n621 34.7936
R5584 avss.n84 avss.n80 34.4123
R5585 avss.n85 avss.n84 34.4123
R5586 avss.n1154 avss.n66 34.4123
R5587 avss.n74 avss.n66 34.4123
R5588 avss.n1240 avss.n1239 34.4123
R5589 avss.n1241 avss.n1240 34.4123
R5590 avss.n38 avss.n37 34.4123
R5591 avss.n1232 avss.n38 34.4123
R5592 avss.n1143 avss.n82 34.4123
R5593 avss.n145 avss.n82 34.4123
R5594 avss.n1139 avss.n90 33.6801
R5595 avss.n1214 avss.t25 33.4847
R5596 avss.t13 avss.n1230 33.4847
R5597 avss.n834 avss.n648 33.1299
R5598 avss.n1211 avss.n48 32.5005
R5599 avss.n1212 avss.n1211 32.5005
R5600 avss.n61 avss.n60 32.5005
R5601 avss.n61 avss.n55 32.5005
R5602 avss.n121 avss.n103 32.5005
R5603 avss.n111 avss.n103 32.5005
R5604 avss.n99 avss.n90 32.5005
R5605 avss.n101 avss.n99 32.5005
R5606 avss.n104 avss.n102 32.5005
R5607 avss.n102 avss.n100 32.5005
R5608 avss.n719 avss.n660 32.0005
R5609 avss.n591 avss.n590 31.6857
R5610 avss.n577 avss.n560 31.6857
R5611 avss.n577 avss.n562 31.6857
R5612 avss.n867 avss.n635 31.2476
R5613 avss.n1247 avss.n1245 30.8082
R5614 avss.n88 avss.n81 30.6755
R5615 avss.n109 avss.n108 30.4899
R5616 avss.n105 avss.n97 30.1319
R5617 avss.n843 avss.n842 30.1181
R5618 avss.n836 avss.n835 30.1181
R5619 avss.n854 avss.n853 30.0632
R5620 avss.n16 avss.n15 29.7851
R5621 avss.n590 avss.n589 29.5874
R5622 avss.n680 avss.n679 29.3652
R5623 avss.n1124 avss.n96 29.3251
R5624 avss.n1075 avss.n168 29.3166
R5625 avss.n621 avss.n604 29.1746
R5626 avss.n707 avss.n706 28.9887
R5627 avss.n705 avss.n704 28.9887
R5628 avss.n843 avss.n643 28.6123
R5629 avss.n828 avss.n650 28.6123
R5630 avss.n1151 avss.n1150 27.7719
R5631 avss.n1152 avss.n1151 27.7719
R5632 avss.n1153 avss.n1152 27.7719
R5633 avss.n1153 avss.n36 27.7719
R5634 avss.n1238 avss.n36 27.7719
R5635 avss.n1238 avss.n1237 27.7719
R5636 avss.n48 avss.n47 26.9228
R5637 avss.n872 avss.n871 26.7299
R5638 avss.n837 avss.n645 26.7299
R5639 avss.n727 avss.n726 25.977
R5640 avss.n147 avss.n140 25.7896
R5641 avss.t57 avss.n1229 25.7367
R5642 avss.n706 avss.n705 25.6005
R5643 avss.n154 avss.n152 25.2546
R5644 avss.n822 avss.n652 24.8476
R5645 avss.n679 avss.n677 24.8476
R5646 avss.n731 avss.n661 24.8476
R5647 avss.n105 avss.n104 24.4927
R5648 avss.n865 avss.n637 24.4711
R5649 avss.n824 avss.n823 24.4711
R5650 avss.n707 avss.n665 24.4711
R5651 avss.n686 avss.n685 24.4711
R5652 avss.n183 avss.n181 24.3755
R5653 avss.n181 avss.n180 24.3755
R5654 avss.n1060 avss.n182 24.3755
R5655 avss.n182 avss.n180 24.3755
R5656 avss.n1129 avss.n1128 24.2648
R5657 avss.n681 avss.n680 24.0946
R5658 avss.n152 avss.n140 23.914
R5659 avss.n842 avss.n841 23.3417
R5660 avss.n855 avss.n854 23.0123
R5661 avss.n861 avss.n637 22.9652
R5662 avss.n823 avss.n822 22.9652
R5663 avss.n915 avss.n914 22.4894
R5664 avss.n914 avss.n184 22.4894
R5665 avss.n1102 avss.n125 22.3548
R5666 avss.n1051 avss.n1022 22.3023
R5667 avss.n140 avss.n139 22.2123
R5668 avss.n867 avss.n866 22.2123
R5669 avss.n147 avss.n30 22.0715
R5670 avss.n1260 avss.n12 22.0326
R5671 avss.n1092 avss.n124 21.7696
R5672 avss.n1102 avss.n126 21.5764
R5673 avss.n22 avss.n21 21.4672
R5674 avss.n16 avss.t6 21.1687
R5675 avss.n1050 avss.n1023 21.1647
R5676 avss.n123 avss.t64 20.9512
R5677 avss.n1036 avss.n1030 20.8934
R5678 avss.n1030 avss.n1029 20.8934
R5679 avss.n837 avss.n836 20.7064
R5680 avss.n786 avss.n785 20.4805
R5681 avss.n785 avss.n765 20.4805
R5682 avss.n773 avss.n765 20.4805
R5683 avss.n731 avss.n660 19.9534
R5684 avss.n608 avss.n233 19.2323
R5685 avss.n630 avss.n629 19.2323
R5686 avss.n847 avss.n643 18.824
R5687 avss.n824 avss.n650 18.824
R5688 avss.n547 avss.n545 18.6433
R5689 avss.n600 avss.n503 18.6433
R5690 avss.n802 avss.n801 18.5384
R5691 avss.n939 avss.n938 18.2862
R5692 avss.n1124 avss.n1123 18.1745
R5693 avss.n835 avss.n834 17.3181
R5694 avss.n47 avss.n43 17.2064
R5695 avss.n1213 avss.n43 17.2064
R5696 avss.n62 avss.n42 17.2064
R5697 avss.n42 avss.n40 17.2064
R5698 avss.n727 avss.n661 16.9417
R5699 avss.t36 avss.n1091 16.8219
R5700 avss.n146 avss.n86 16.2505
R5701 avss.n146 avss.t41 16.2505
R5702 avss.n143 avss.n142 16.2505
R5703 avss.t41 avss.n143 16.2505
R5704 avss.n22 avss.n15 16.1338
R5705 avss.n1110 avss.n120 16.0005
R5706 avss.n1117 avss.n97 15.7807
R5707 avss.n1135 avss.n1124 15.7807
R5708 avss.n1088 avss.n159 15.5506
R5709 avss.n1116 avss.n1115 15.4875
R5710 avss.n1221 avss.n1220 15.4479
R5711 avss.n873 avss.n872 15.4358
R5712 avss.n155 avss.n154 15.3345
R5713 avss.n1115 avss.n1114 15.0967
R5714 avss.n548 avss.n508 15.0005
R5715 avss.n508 avss.n506 15.0005
R5716 avss.n510 avss.n507 15.0005
R5717 avss.n507 avss.n506 15.0005
R5718 avss.n504 avss.n501 15.0005
R5719 avss.n582 avss.n501 15.0005
R5720 avss.n599 avss.n502 15.0005
R5721 avss.n582 avss.n502 15.0005
R5722 avss.n1040 avss.n1023 14.7701
R5723 avss.n687 avss.n686 14.6829
R5724 avss.n76 avss.n32 14.6255
R5725 avss.n77 avss.n76 14.6255
R5726 avss.n1159 avss.n1158 14.6255
R5727 avss.n1160 avss.n1159 14.6255
R5728 avss.n523 avss.n519 14.5302
R5729 avss.n206 avss.n205 14.448
R5730 avss.n925 avss.n198 14.3554
R5731 avss.n830 avss.n648 14.3064
R5732 avss.n631 avss.n630 14.1378
R5733 avss.n801 avss.n800 13.9481
R5734 avss.n800 avss.n738 13.9481
R5735 avss.n759 avss.n738 13.9481
R5736 avss.n760 avss.n759 13.9481
R5737 avss.n787 avss.n786 13.9481
R5738 avss.n1093 avss.n126 13.6799
R5739 avss.n1254 avss.n1253 13.6052
R5740 avss.n1255 avss.n1254 13.6052
R5741 avss.n144 avss.n79 13.6052
R5742 avss.n144 avss.n73 13.6052
R5743 avss.n1244 avss.n1243 13.6052
R5744 avss.n1243 avss.n1242 13.6052
R5745 avss.n148 avss.n147 13.6052
R5746 avss.n149 avss.n148 13.6052
R5747 avss.n174 avss.n169 13.6052
R5748 avss.n174 avss.n173 13.6052
R5749 avss.n170 avss.n168 13.6052
R5750 avss.n173 avss.n170 13.6052
R5751 avss.n1084 avss.n162 13.6052
R5752 avss.n164 avss.n161 13.6052
R5753 avss.n1080 avss.n161 13.6052
R5754 avss.n608 avss.n605 13.5647
R5755 avss.n52 avss.n51 13.5534
R5756 avss.n518 avss.n514 13.2848
R5757 avss.n1081 avss.n162 13.0635
R5758 avss.n694 avss.n670 12.424
R5759 avss.n51 avss.n11 12.1845
R5760 avss.n1261 avss.n11 12.0414
R5761 avss.n1114 avss.n113 11.9211
R5762 avss.t69 avss.t16 11.5374
R5763 avss.n1260 avss.n1259 11.4592
R5764 avss.n60 avss.n3 11.405
R5765 avss.n718 avss.n717 11.2946
R5766 avss.n829 avss.n828 11.2946
R5767 avss.n713 avss.n712 11.2946
R5768 avss.n1245 avss.n31 11.2477
R5769 avss.n1040 avss.n1039 11.2225
R5770 avss.n141 avss.n31 10.912
R5771 avss.n1135 avss.n1134 10.6509
R5772 avss.n1134 avss.n1133 10.6509
R5773 avss.n1123 avss.n97 10.4066
R5774 avss.n1092 avss.n113 10.26
R5775 avss.n47 avss.n45 10.1559
R5776 avss.n933 avss.n194 9.75892
R5777 avss.n1230 avss.t24 9.74291
R5778 avss.n1214 avss.t17 9.74291
R5779 avss.n522 avss.n193 9.63218
R5780 avss.n28 avss.n26 9.59066
R5781 avss.t34 avss.n26 9.59066
R5782 avss.n1246 avss.n25 9.59066
R5783 avss.t34 avss.n25 9.59066
R5784 avss.n1038 avss.n1022 9.35596
R5785 dvss avss.n677 9.3308
R5786 avss.n410 avss.n264 9.30106
R5787 avss.n453 avss.n243 9.30106
R5788 avss.n387 avss.n276 9.30106
R5789 avss.n362 avss.n313 9.30106
R5790 avss.n480 avss.n479 9.30101
R5791 avss.n340 avss.n339 9.30101
R5792 avss.n726 avss.n725 9.3005
R5793 avss.n679 avss.n678 9.3005
R5794 avss.n680 avss.n676 9.3005
R5795 avss.n682 avss.n681 9.3005
R5796 avss.n683 avss.n675 9.3005
R5797 avss.n685 avss.n684 9.3005
R5798 avss.n686 avss.n674 9.3005
R5799 avss.n687 avss.n673 9.3005
R5800 avss.n689 avss.n688 9.3005
R5801 avss.n690 avss.n672 9.3005
R5802 avss.n692 avss.n691 9.3005
R5803 avss.n693 avss.n671 9.3005
R5804 avss.n695 avss.n694 9.3005
R5805 avss.n696 avss.n670 9.3005
R5806 avss.n698 avss.n697 9.3005
R5807 avss.n699 avss.n669 9.3005
R5808 avss.n701 avss.n700 9.3005
R5809 avss.n702 avss.n668 9.3005
R5810 avss.n704 avss.n703 9.3005
R5811 avss.n705 avss.n667 9.3005
R5812 avss.n706 avss.n666 9.3005
R5813 avss.n708 avss.n707 9.3005
R5814 avss.n709 avss.n665 9.3005
R5815 avss.n711 avss.n710 9.3005
R5816 avss.n712 avss.n664 9.3005
R5817 avss.n714 avss.n713 9.3005
R5818 avss.n715 avss.n663 9.3005
R5819 avss.n717 avss.n716 9.3005
R5820 avss.n718 avss.n662 9.3005
R5821 avss.n720 avss.n719 9.3005
R5822 avss.n729 avss.n661 9.3005
R5823 avss.n728 avss.n727 9.3005
R5824 avss.n726 avss.n722 9.3005
R5825 avss.n731 avss.n730 9.3005
R5826 avss.n288 avss.n287 9.3005
R5827 avss.n287 avss.n286 9.3005
R5828 avss.n287 avss.n284 9.3005
R5829 avss.n299 avss.n298 9.3005
R5830 avss.n298 avss.n297 9.3005
R5831 avss.n298 avss.n296 9.3005
R5832 avss.n310 avss.n309 9.3005
R5833 avss.n309 avss.n308 9.3005
R5834 avss.n309 avss.n307 9.3005
R5835 avss.n325 avss.n324 9.3005
R5836 avss.n324 avss.n323 9.3005
R5837 avss.n324 avss.n322 9.3005
R5838 avss.n336 avss.n335 9.3005
R5839 avss.n335 avss.n334 9.3005
R5840 avss.n335 avss.n332 9.3005
R5841 avss.n394 avss.n393 9.3005
R5842 avss.n272 avss.n271 9.3005
R5843 avss.n386 avss.n277 9.3005
R5844 avss.n385 avss.n278 9.3005
R5845 avss.n285 avss.n279 9.3005
R5846 avss.n379 avss.n283 9.3005
R5847 avss.n378 avss.n289 9.3005
R5848 avss.n377 avss.n290 9.3005
R5849 avss.n295 avss.n291 9.3005
R5850 avss.n371 avss.n300 9.3005
R5851 avss.n370 avss.n301 9.3005
R5852 avss.n369 avss.n302 9.3005
R5853 avss.n311 avss.n303 9.3005
R5854 avss.n363 avss.n312 9.3005
R5855 avss.n361 avss.n314 9.3005
R5856 avss.n321 avss.n315 9.3005
R5857 avss.n355 avss.n319 9.3005
R5858 avss.n354 avss.n320 9.3005
R5859 avss.n353 avss.n326 9.3005
R5860 avss.n333 avss.n327 9.3005
R5861 avss.n347 avss.n331 9.3005
R5862 avss.n346 avss.n337 9.3005
R5863 avss.n345 avss.n338 9.3005
R5864 avss.n425 avss.n424 9.3005
R5865 avss.n424 avss.n423 9.3005
R5866 avss.n424 avss.n259 9.3005
R5867 avss.n429 avss.n252 9.3005
R5868 avss.n430 avss.n429 9.3005
R5869 avss.n429 avss.n427 9.3005
R5870 avss.n443 avss.n442 9.3005
R5871 avss.n442 avss.n251 9.3005
R5872 avss.n442 avss.n441 9.3005
R5873 avss.n492 avss.n491 9.3005
R5874 avss.n492 avss.n455 9.3005
R5875 avss.n493 avss.n492 9.3005
R5876 avss.n485 avss.n484 9.3005
R5877 avss.n486 avss.n485 9.3005
R5878 avss.n485 avss.n457 9.3005
R5879 avss.n266 avss.n265 9.3005
R5880 avss.n409 avss.n408 9.3005
R5881 avss.n413 avss.n412 9.3005
R5882 avss.n411 avss.n260 9.3005
R5883 avss.n422 avss.n421 9.3005
R5884 avss.n420 avss.n258 9.3005
R5885 avss.n426 avss.n257 9.3005
R5886 avss.n432 avss.n431 9.3005
R5887 avss.n428 avss.n253 9.3005
R5888 avss.n439 avss.n438 9.3005
R5889 avss.n440 avss.n250 9.3005
R5890 avss.n445 avss.n444 9.3005
R5891 avss.n246 avss.n245 9.3005
R5892 avss.n452 avss.n451 9.3005
R5893 avss.n496 avss.n495 9.3005
R5894 avss.n494 avss.n244 9.3005
R5895 avss.n467 avss.n454 9.3005
R5896 avss.n458 avss.n456 9.3005
R5897 avss.n490 avss.n489 9.3005
R5898 avss.n488 avss.n487 9.3005
R5899 avss.n462 avss.n461 9.3005
R5900 avss.n483 avss.n482 9.3005
R5901 avss.n481 avss.n463 9.3005
R5902 avss.n820 avss.n652 9.3005
R5903 avss.n874 avss.n873 9.3005
R5904 avss.n872 avss.n634 9.3005
R5905 avss.n871 avss.n870 9.3005
R5906 avss.n869 avss.n635 9.3005
R5907 avss.n868 avss.n867 9.3005
R5908 avss.n866 avss.n636 9.3005
R5909 avss.n865 avss.n864 9.3005
R5910 avss.n863 avss.n637 9.3005
R5911 avss.n862 avss.n861 9.3005
R5912 avss.n860 avss.n638 9.3005
R5913 avss.n859 avss.n858 9.3005
R5914 avss.n857 avss.n639 9.3005
R5915 avss.n856 avss.n855 9.3005
R5916 avss.n854 avss.n640 9.3005
R5917 avss.n853 avss.n852 9.3005
R5918 avss.n851 avss.n641 9.3005
R5919 avss.n850 avss.n849 9.3005
R5920 avss.n848 avss.n642 9.3005
R5921 avss.n847 avss.n846 9.3005
R5922 avss.n845 avss.n643 9.3005
R5923 avss.n844 avss.n843 9.3005
R5924 avss.n842 avss.n644 9.3005
R5925 avss.n841 avss.n840 9.3005
R5926 avss.n839 avss.n645 9.3005
R5927 avss.n838 avss.n837 9.3005
R5928 avss.n836 avss.n646 9.3005
R5929 avss.n835 avss.n647 9.3005
R5930 avss.n834 avss.n833 9.3005
R5931 avss.n832 avss.n648 9.3005
R5932 avss.n831 avss.n830 9.3005
R5933 avss.n829 avss.n649 9.3005
R5934 avss.n828 avss.n827 9.3005
R5935 avss.n826 avss.n650 9.3005
R5936 avss.n825 avss.n824 9.3005
R5937 avss.n823 avss.n651 9.3005
R5938 avss.n822 avss.n821 9.3005
R5939 avss.n885 avss.n226 8.79354
R5940 avss.n1138 avss.n88 8.58924
R5941 avss.n922 avss.n921 8.19036
R5942 avss.n212 avss.n211 8.18274
R5943 avss.n929 avss.n199 8.18274
R5944 avss.n1093 avss.n1092 8.15928
R5945 avss.n132 avss.n126 8.11042
R5946 avss.n1139 avss.n1138 8.03513
R5947 avss.n1076 avss.n167 7.82362
R5948 avss.n762 avss.n760 7.6805
R5949 avss.n1106 avss.n112 7.49854
R5950 avss.n1110 avss.n1109 7.34571
R5951 avss.n1074 avss.n1073 7.13465
R5952 avss.n172 avss.n171 7.13465
R5953 avss.n172 avss.n160 7.13465
R5954 avss.n1086 avss.n1085 7.13465
R5955 avss.n1087 avss.n1086 7.13465
R5956 avss.n1083 avss.n1082 7.13465
R5957 avss.n1128 avss.n88 7.01267
R5958 avss.n58 avss.n11 6.69588
R5959 avss.n96 avss.n90 6.4005
R5960 avss.n1036 avss.n1031 6.28553
R5961 avss.n787 avss.n762 6.26809
R5962 avss.n395 avss.n270 6.13547
R5963 avss.n401 avss.n400 6.13534
R5964 avss.n878 avss.n226 5.89963
R5965 avss.n59 avss.n58 5.61281
R5966 avss.n598 avss.n596 5.6005
R5967 avss.n1042 avss.n1041 5.51906
R5968 avss.n549 avss.n509 5.4005
R5969 avss.t60 avss.n145 5.32523
R5970 avss.n85 avss.t33 5.32523
R5971 avss.n1027 avss.n1025 5.13208
R5972 avss.n1045 avss.n1027 5.13208
R5973 avss.n631 avss.n233 5.09503
R5974 avss.n1103 avss.n1102 5.08147
R5975 avss.n934 avss.n193 5.06981
R5976 avss.n1147 avss.n1145 5.05494
R5977 avss.n1234 avss.n1233 5.02119
R5978 avss.n934 avss.n933 4.94307
R5979 avss.n1103 avss.n124 4.86695
R5980 avss.n1227 avss.n44 4.66041
R5981 avss.n1039 avss.n1038 4.65428
R5982 avss.n721 avss.n660 4.6359
R5983 avss.n1147 avss.n1146 4.46947
R5984 avss.n1234 avss.n35 4.46947
R5985 avss.n598 avss.n597 4.38075
R5986 avss.n546 avss.n509 4.37879
R5987 avss.n18 avss.n13 4.36669
R5988 avss.n123 avss.n122 4.36128
R5989 avss.n1146 avss.n68 4.30062
R5990 avss.n1021 avss.n1019 4.29698
R5991 avss.n1037 avss.n1035 4.21607
R5992 avss.n1035 avss.n1034 4.14944
R5993 avss.n1034 avss.n1033 4.14944
R5994 avss.n1026 avss.n1024 4.09141
R5995 avss.n1028 avss.n1026 4.09141
R5996 avss.n523 avss.n522 3.91448
R5997 avss.n1059 avss.n184 3.91161
R5998 avss.n1248 avss.n30 3.67161
R5999 avss.n1157 avss.n1156 3.66244
R6000 avss.n1231 avss.t43 3.55032
R6001 avss.n1259 avss.n13 3.50683
R6002 avss.n1032 avss.n1024 3.34378
R6003 avss.n818 avss.n817 3.27492
R6004 avss.n1129 avss.n81 3.22833
R6005 avss.n1165 avss.n1164 3.05772
R6006 avss.n65 avss.n35 3.05584
R6007 avss.n1077 avss.n1076 2.98691
R6008 avss.n1251 avss.n29 2.94732
R6009 avss.n1249 avss.n1248 2.91148
R6010 avss.n879 avss.n878 2.89441
R6011 avss.n121 avss.n112 2.87229
R6012 avss.n60 avss.n59 2.86873
R6013 avss.n21 avss.n20 2.80414
R6014 avss.n1144 avss.n1143 2.61868
R6015 avss.n587 avss.n232 2.60526
R6016 avss.n1142 avss.n1141 2.47323
R6017 avss.n1141 avss.n88 2.47323
R6018 avss.n122 avss.n112 2.44756
R6019 avss.n588 avss.n558 2.35044
R6020 avss.n633 avss.n231 2.19136
R6021 avss.n586 avss.n585 2.17408
R6022 avss.n1058 avss.n940 2.15152
R6023 avss.n1108 avss.n120 2.1169
R6024 avss.n589 avss.n560 2.09886
R6025 avss.n49 avss.n12 2.05207
R6026 avss.n63 avss.n29 1.93399
R6027 avss.n107 avss.n104 1.89703
R6028 avss.n108 avss.n107 1.89382
R6029 avss.n819 avss.n818 1.8605
R6030 avss.n1107 avss.n1106 1.8605
R6031 avss.n106 avss.n105 1.8605
R6032 avss.n1117 avss.n1116 1.85699
R6033 avss.n1021 avss.n1020 1.82489
R6034 avss.n1058 avss.n1057 1.81171
R6035 avss.n1251 avss.n1250 1.72169
R6036 avss.n400 avss.n265 1.64187
R6037 avss.n395 avss.n394 1.64057
R6038 avss.n1077 avss.n165 1.5837
R6039 avss.n1043 avss.n1042 1.56886
R6040 avss.n1044 avss.n1043 1.56886
R6041 avss.n1206 avss.n1205 1.5505
R6042 avss.n1266 avss.n4 1.49704
R6043 avss.n546 avss.n231 1.49237
R6044 avss avss.n1 1.48104
R6045 avss.n875 avss.n874 1.45077
R6046 avss.n569 avss.n558 1.44956
R6047 dvss avss.n230 1.44157
R6048 avss.n1225 avss.n1224 1.32133
R6049 avss.n1270 avss.n1269 1.31102
R6050 avss.n761 avss.n653 1.30418
R6051 avss.n876 avss.n230 1.29478
R6052 avss.n1104 avss.n123 1.28462
R6053 avss.n519 avss.n518 1.24591
R6054 avss.n1167 avss 1.23982
R6055 avss.n587 avss.n586 1.23022
R6056 avss.n588 avss.n587 1.22373
R6057 avss.n518 avss.n517 1.22095
R6058 avss.n1049 avss.n1048 1.20521
R6059 avss.n1203 avss.n1202 1.19172
R6060 avss.n597 avss.n232 1.15531
R6061 avss.n1048 avss.n1047 1.13422
R6062 avss.n1047 avss.n1046 1.13422
R6063 avss.n1164 avss.n65 1.09236
R6064 avss.n1266 avss.n1265 1.06941
R6065 avss.n819 avss.n653 1.0534
R6066 avss.n878 avss.n877 1.01717
R6067 avss.n20 avss.n19 0.957122
R6068 avss.n167 avss.n166 0.936734
R6069 avss.n1158 avss.n79 0.893523
R6070 avss.n819 dvss 0.86713
R6071 avss.n17 avss.n16 0.845955
R6072 avss.n46 avss.n44 0.845955
R6073 avss.n1244 avss.n32 0.841376
R6074 avss.n999 avss.n998 0.837244
R6075 avss.n1052 avss.n1021 0.808157
R6076 dvss avss.n653 0.733375
R6077 avss.n1168 avss.n62 0.731929
R6078 avss.n164 avss.n163 0.714663
R6079 dvss avss.n230 0.71054
R6080 avss.n1225 avss.n46 0.686469
R6081 avss.n1056 avss.n1054 0.681951
R6082 avss.n1057 dvss 0.679512
R6083 avss.n1155 avss.n64 0.672416
R6084 avss.n1220 avss.n3 0.650441
R6085 avss.n1250 avss.n1249 0.634111
R6086 avss.n1057 avss.n1056 0.626581
R6087 avss.n1226 avss.n1225 0.6205
R6088 avss.n17 avss.n4 0.606103
R6089 avss.n1169 avss.n1167 0.604749
R6090 avss.n940 avss.n939 0.603757
R6091 avss.n632 avss.n631 0.603227
R6092 avss.n1267 avss.n3 0.593683
R6093 avss.n1053 avss.n167 0.584781
R6094 avss.n1202 avss.n1201 0.582318
R6095 avss.n1269 avss 0.566822
R6096 avss.n1053 avss.n1052 0.53923
R6097 avss.n1056 avss.n1055 0.539165
R6098 avss.n1081 avss.n1080 0.536142
R6099 avss.n1224 avss.n1223 0.517167
R6100 avss.n1109 avss.n1108 0.517167
R6101 avss.n517 avss.n516 0.516217
R6102 avss.n1150 avss.n81 0.457643
R6103 avss.n1019 avss.n1018 0.450328
R6104 avss.n998 avss.n978 0.438865
R6105 avss.n1109 avss.n121 0.438107
R6106 avss.n1076 avss.n1075 0.407877
R6107 avss.n1205 avss.n1169 0.406136
R6108 avss.n589 avss.n588 0.404848
R6109 avss.n1204 avss.n1203 0.398755
R6110 avss.n1224 avss.n2 0.39776
R6111 avss.n940 avss.n185 0.396762
R6112 avss.n19 avss.n18 0.389389
R6113 avss.n1204 avss.n2 0.388725
R6114 avss.n1157 avss.n68 0.386852
R6115 avss.n1156 avss.n63 0.358192
R6116 dvss avss.n819 0.356294
R6117 avss.n1165 avss.n64 0.353256
R6118 avss.n1039 avss.n1031 0.344944
R6119 avss.n1107 avss.n1105 0.335899
R6120 avss.n106 avss.n1 0.32778
R6121 avss.n107 avss.n106 0.323689
R6122 avss.n1166 avss.n1165 0.3105
R6123 avss.n1169 avss.n1168 0.3005
R6124 avss.n762 avss.n761 0.3005
R6125 avss.n153 avss.n29 0.298417
R6126 avss.n1104 avss.n1103 0.293439
R6127 avss.n877 dvss 0.2894
R6128 avss.n1108 avss.n1107 0.288899
R6129 avss.n1059 avss.n1058 0.284911
R6130 avss.n1268 avss.n2 0.28415
R6131 avss.n1078 avss.n164 0.275178
R6132 avss.n517 avss.n185 0.272299
R6133 avss.n1252 avss.n1251 0.266214
R6134 avss.n1203 avss 0.260623
R6135 avss.n18 avss.n17 0.256966
R6136 avss.n205 avss.n194 0.253965
R6137 avss.n206 avss.n198 0.253965
R6138 avss.n548 avss.n547 0.238561
R6139 avss.n504 avss.n503 0.238561
R6140 avss.n1078 avss.n1077 0.221929
R6141 avss.n1250 avss.n27 0.207167
R6142 avss.n1167 avss.n46 0.20273
R6143 avss.n1116 avss.n0 0.179346
R6144 avss avss.n1266 0.173899
R6145 avss.n877 avss.n876 0.170624
R6146 avss.n1253 avss.n27 0.163557
R6147 avss.n516 avss.n231 0.16209
R6148 avss.n1270 avss.n1 0.152695
R6149 avss.n875 avss.n633 0.149407
R6150 avss.n1105 avss.n1104 0.148401
R6151 avss.n761 avss.n165 0.129071
R6152 avss.n876 avss.n875 0.119023
R6153 dvss avss.n1053 0.118752
R6154 avss.n1170 avss 0.114272
R6155 avss.n1205 avss.n1204 0.109693
R6156 avss.n1223 avss.n48 0.106285
R6157 avss.n943 avss.n941 0.10275
R6158 avss.n962 avss.n960 0.10275
R6159 avss.n981 avss.n979 0.10275
R6160 avss.n1002 avss.n1000 0.10275
R6161 avss.n165 dvss 0.0930926
R6162 avss.n721 avss.n720 0.0918107
R6163 avss.n1025 avss.n1023 0.0907913
R6164 avss.n1267 avss 0.0896768
R6165 avss.n1248 avss.n1247 0.0866111
R6166 dvss avss.n185 0.084875
R6167 avss.n632 avss.n232 0.0835912
R6168 avss.n998 avss.n997 0.0788906
R6169 avss.n633 avss.n632 0.0765474
R6170 avss.n1105 avss.n0 0.0758817
R6171 avss.n516 dvss 0.0731595
R6172 avss.n1038 avss.n1037 0.0709545
R6173 avss.n1032 avss.n1022 0.0704248
R6174 avss.n945 avss.n943 0.06865
R6175 avss.n947 avss.n945 0.06865
R6176 avss.n949 avss.n947 0.06865
R6177 avss.n951 avss.n949 0.06865
R6178 avss.n953 avss.n951 0.06865
R6179 avss.n955 avss.n953 0.06865
R6180 avss.n957 avss.n955 0.06865
R6181 avss.n959 avss.n957 0.06865
R6182 avss.n964 avss.n962 0.06865
R6183 avss.n966 avss.n964 0.06865
R6184 avss.n968 avss.n966 0.06865
R6185 avss.n970 avss.n968 0.06865
R6186 avss.n972 avss.n970 0.06865
R6187 avss.n974 avss.n972 0.06865
R6188 avss.n976 avss.n974 0.06865
R6189 avss.n978 avss.n976 0.06865
R6190 avss.n983 avss.n981 0.06865
R6191 avss.n985 avss.n983 0.06865
R6192 avss.n987 avss.n985 0.06865
R6193 avss.n989 avss.n987 0.06865
R6194 avss.n991 avss.n989 0.06865
R6195 avss.n993 avss.n991 0.06865
R6196 avss.n995 avss.n993 0.06865
R6197 avss.n997 avss.n995 0.06865
R6198 avss.n1004 avss.n1002 0.06865
R6199 avss.n1006 avss.n1004 0.06865
R6200 avss.n1008 avss.n1006 0.06865
R6201 avss.n1010 avss.n1008 0.06865
R6202 avss.n1012 avss.n1010 0.06865
R6203 avss.n1014 avss.n1012 0.06865
R6204 avss.n1016 avss.n1014 0.06865
R6205 avss.n1018 avss.n1016 0.06865
R6206 avss.n999 avss.n959 0.0632125
R6207 dvss avss.n721 0.0615076
R6208 avss.n678 avss.n676 0.0611061
R6209 avss.n682 avss.n676 0.0611061
R6210 avss.n683 avss.n682 0.0611061
R6211 avss.n684 avss.n683 0.0611061
R6212 avss.n684 avss.n674 0.0611061
R6213 avss.n674 avss.n673 0.0611061
R6214 avss.n689 avss.n673 0.0611061
R6215 avss.n690 avss.n689 0.0611061
R6216 avss.n691 avss.n690 0.0611061
R6217 avss.n691 avss.n671 0.0611061
R6218 avss.n695 avss.n671 0.0611061
R6219 avss.n696 avss.n695 0.0611061
R6220 avss.n697 avss.n696 0.0611061
R6221 avss.n697 avss.n669 0.0611061
R6222 avss.n701 avss.n669 0.0611061
R6223 avss.n702 avss.n701 0.0611061
R6224 avss.n703 avss.n702 0.0611061
R6225 avss.n703 avss.n667 0.0611061
R6226 avss.n667 avss.n666 0.0611061
R6227 avss.n708 avss.n666 0.0611061
R6228 avss.n709 avss.n708 0.0611061
R6229 avss.n710 avss.n709 0.0611061
R6230 avss.n714 avss.n664 0.0611061
R6231 avss.n715 avss.n714 0.0611061
R6232 avss.n716 avss.n715 0.0611061
R6233 avss.n716 avss.n662 0.0611061
R6234 avss.n720 avss.n662 0.0611061
R6235 avss.n729 avss.n728 0.0611061
R6236 avss.n728 avss.n722 0.0611061
R6237 avss.n870 avss.n634 0.0550455
R6238 avss.n870 avss.n869 0.0550455
R6239 avss.n869 avss.n868 0.0550455
R6240 avss.n868 avss.n636 0.0550455
R6241 avss.n864 avss.n636 0.0550455
R6242 avss.n864 avss.n863 0.0550455
R6243 avss.n863 avss.n862 0.0550455
R6244 avss.n862 avss.n638 0.0550455
R6245 avss.n858 avss.n638 0.0550455
R6246 avss.n858 avss.n857 0.0550455
R6247 avss.n857 avss.n856 0.0550455
R6248 avss.n856 avss.n640 0.0550455
R6249 avss.n852 avss.n640 0.0550455
R6250 avss.n852 avss.n851 0.0550455
R6251 avss.n851 avss.n850 0.0550455
R6252 avss.n850 avss.n642 0.0550455
R6253 avss.n846 avss.n642 0.0550455
R6254 avss.n846 avss.n845 0.0550455
R6255 avss.n845 avss.n844 0.0550455
R6256 avss.n844 avss.n644 0.0550455
R6257 avss.n840 avss.n644 0.0550455
R6258 avss.n840 avss.n839 0.0550455
R6259 avss.n838 avss.n646 0.0550455
R6260 avss.n647 avss.n646 0.0550455
R6261 avss.n833 avss.n647 0.0550455
R6262 avss.n833 avss.n832 0.0550455
R6263 avss.n832 avss.n831 0.0550455
R6264 avss.n831 avss.n649 0.0550455
R6265 avss.n827 avss.n649 0.0550455
R6266 avss.n827 avss.n826 0.0550455
R6267 avss.n826 avss.n825 0.0550455
R6268 avss.n825 avss.n651 0.0550455
R6269 avss.n821 avss.n651 0.0550455
R6270 avss.n412 avss.n410 0.0546569
R6271 avss.n495 avss.n453 0.0546569
R6272 avss.n479 avss.n463 0.0537932
R6273 avss.n410 avss.n409 0.0537291
R6274 avss.n453 avss.n452 0.0537291
R6275 avss.n277 avss.n276 0.0535264
R6276 avss.n314 avss.n313 0.0535264
R6277 avss.n409 avss.n265 0.0533634
R6278 avss.n412 avss.n411 0.0533634
R6279 avss.n440 avss.n439 0.0533634
R6280 avss.n452 avss.n245 0.0533634
R6281 avss.n495 avss.n494 0.0533634
R6282 avss.n483 avss.n463 0.0533634
R6283 avss.n339 avss.n338 0.0526569
R6284 avss.n276 avss.n271 0.0525955
R6285 avss.n313 avss.n312 0.0525955
R6286 avss.n394 avss.n271 0.0522241
R6287 avss.n278 avss.n277 0.0522241
R6288 avss.n301 avss.n300 0.0522241
R6289 avss.n312 avss.n311 0.0522241
R6290 avss.n321 avss.n314 0.0522241
R6291 avss.n338 avss.n337 0.0522241
R6292 avss.n724 dvss 0.0503737
R6293 avss avss.n1166 0.0500072
R6294 avss.n427 avss.n426 0.0484075
R6295 avss.n490 avss.n457 0.0484075
R6296 avss.n296 avss.n289 0.047375
R6297 avss.n332 avss.n326 0.047375
R6298 avss.n426 avss.n425 0.0451035
R6299 avss.n491 avss.n490 0.0451035
R6300 avss.n289 avss.n288 0.0441422
R6301 avss.n326 avss.n325 0.0441422
R6302 avss.n1269 avss.n1268 0.0421667
R6303 avss.n724 avss.n722 0.0415354
R6304 avss.n1052 avss.n1051 0.0392931
R6305 avss.n411 avss.n259 0.0351916
R6306 avss.n431 avss.n430 0.0351916
R6307 avss.n444 avss.n443 0.0351916
R6308 avss.n494 avss.n493 0.0351916
R6309 avss.n487 avss.n486 0.0351916
R6310 avss.n943 avss.n942 0.0346
R6311 avss.n945 avss.n944 0.0346
R6312 avss.n947 avss.n946 0.0346
R6313 avss.n949 avss.n948 0.0346
R6314 avss.n951 avss.n950 0.0346
R6315 avss.n953 avss.n952 0.0346
R6316 avss.n955 avss.n954 0.0346
R6317 avss.n957 avss.n956 0.0346
R6318 avss.n959 avss.n958 0.0346
R6319 avss.n962 avss.n961 0.0346
R6320 avss.n964 avss.n963 0.0346
R6321 avss.n966 avss.n965 0.0346
R6322 avss.n968 avss.n967 0.0346
R6323 avss.n970 avss.n969 0.0346
R6324 avss.n972 avss.n971 0.0346
R6325 avss.n974 avss.n973 0.0346
R6326 avss.n976 avss.n975 0.0346
R6327 avss.n978 avss.n977 0.0346
R6328 avss.n981 avss.n980 0.0346
R6329 avss.n983 avss.n982 0.0346
R6330 avss.n985 avss.n984 0.0346
R6331 avss.n987 avss.n986 0.0346
R6332 avss.n989 avss.n988 0.0346
R6333 avss.n991 avss.n990 0.0346
R6334 avss.n993 avss.n992 0.0346
R6335 avss.n995 avss.n994 0.0346
R6336 avss.n997 avss.n996 0.0346
R6337 avss.n1002 avss.n1001 0.0346
R6338 avss.n1004 avss.n1003 0.0346
R6339 avss.n1006 avss.n1005 0.0346
R6340 avss.n1008 avss.n1007 0.0346
R6341 avss.n1010 avss.n1009 0.0346
R6342 avss.n1012 avss.n1011 0.0346
R6343 avss.n1014 avss.n1013 0.0346
R6344 avss.n1016 avss.n1015 0.0346
R6345 avss.n1018 avss.n1017 0.0346
R6346 avss.n284 avss.n278 0.034444
R6347 avss.n297 avss.n290 0.034444
R6348 avss.n310 avss.n302 0.034444
R6349 avss.n322 avss.n321 0.034444
R6350 avss.n334 avss.n333 0.034444
R6351 avss.n1156 avss.n1155 0.0340958
R6352 avss.n423 avss.n258 0.0318877
R6353 avss.n439 avss.n252 0.0318877
R6354 avss.n456 avss.n455 0.0318877
R6355 avss.n484 avss.n483 0.0318877
R6356 avss avss.n1170 0.03175
R6357 avss.n286 avss.n283 0.0312112
R6358 avss.n300 avss.n299 0.0312112
R6359 avss.n323 avss.n320 0.0312112
R6360 avss.n337 avss.n336 0.0312112
R6361 avss.n678 dvss 0.030803
R6362 avss.n710 dvss 0.030803
R6363 dvss avss.n664 0.030803
R6364 avss.n730 dvss 0.030803
R6365 avss.n730 dvss 0.030803
R6366 dvss avss.n729 0.030803
R6367 avss.n874 dvss 0.0277727
R6368 avss.n634 dvss 0.0277727
R6369 avss.n839 dvss 0.0277727
R6370 dvss avss.n838 0.0277727
R6371 avss.n821 dvss 0.0277727
R6372 dvss avss.n820 0.0277727
R6373 avss.n820 dvss 0.0277727
R6374 avss.n479 dvss 0.0274177
R6375 avss.n339 dvss 0.0268486
R6376 avss.n1041 avss.n1040 0.0266972
R6377 avss.n725 dvss 0.0246935
R6378 avss.n423 avss.n422 0.0219758
R6379 avss.n428 avss.n252 0.0219758
R6380 dvss avss.n251 0.0219758
R6381 avss.n455 avss.n454 0.0219758
R6382 avss.n484 avss.n462 0.0219758
R6383 avss.n286 avss.n285 0.0215129
R6384 avss.n299 avss.n295 0.0215129
R6385 avss.n308 dvss 0.0215129
R6386 avss.n323 avss.n319 0.0215129
R6387 avss.n336 avss.n331 0.0215129
R6388 avss.n1050 avss.n1049 0.0196358
R6389 avss.n422 avss.n259 0.0186718
R6390 avss.n430 avss.n428 0.0186718
R6391 avss.n441 dvss 0.0186718
R6392 avss.n443 avss.n245 0.0186718
R6393 avss.n493 avss.n454 0.0186718
R6394 avss.n486 avss.n462 0.0186718
R6395 avss.n285 avss.n284 0.0182802
R6396 avss.n297 avss.n295 0.0182802
R6397 dvss avss.n307 0.0182802
R6398 avss.n311 avss.n310 0.0182802
R6399 avss.n322 avss.n319 0.0182802
R6400 avss.n334 avss.n331 0.0182802
R6401 avss.n1268 avss.n1267 0.0176494
R6402 avss.n725 avss.n724 0.016125
R6403 avss.n1166 avss.n63 0.0146129
R6404 avss avss.n0 0.0133817
R6405 avss.n547 avss.n546 0.0125063
R6406 avss.n597 avss.n503 0.0125063
R6407 avss avss.n1270 0.0119504
R6408 avss.n19 avss.n4 0.00875991
R6409 avss.n425 avss.n258 0.00875991
R6410 avss.n441 avss.n440 0.00875991
R6411 avss.n491 avss.n456 0.00875991
R6412 avss.n288 avss.n283 0.0085819
R6413 avss.n307 avss.n301 0.0085819
R6414 avss.n325 avss.n320 0.0085819
R6415 avss.n1051 avss.n1050 0.00626923
R6416 avss.n431 avss.n427 0.00545595
R6417 avss.n444 avss.n251 0.00545595
R6418 avss.n487 avss.n457 0.00545595
R6419 avss.n296 avss.n290 0.00534914
R6420 avss.n308 avss.n302 0.00534914
R6421 avss.n333 avss.n332 0.00534914
R6422 avss.n1019 avss.n999 0.00291667
R6423 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n47 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n46 156.462
R6424 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n54 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n53 156.462
R6425 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n38 69.6745
R6426 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n1 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n4 69.6745
R6427 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n41 69.6745
R6428 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n0 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n42 69.6745
R6429 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n37 69.6745
R6430 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n12 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A 69.6745
R6431 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n1 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n36 69.6745
R6432 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n7 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n1 69.6745
R6433 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n40 69.6745
R6434 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n27 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A 69.6745
R6435 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n0 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n39 69.6745
R6436 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n22 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n0 69.6745
R6437 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n48 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n44 155.492
R6438 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n55 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n51 155.492
R6439 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n45 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t33 113.543
R6440 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n52 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t47 113.543
R6441 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n50 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t60 93.5093
R6442 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n43 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t46 93.5085
R6443 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n2 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t32 92.5445
R6444 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n3 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t55 92.5445
R6445 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n5 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t30 92.5445
R6446 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n6 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t54 92.5445
R6447 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n8 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t4 92.5445
R6448 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n9 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t31 92.5445
R6449 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n10 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t38 92.5445
R6450 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n11 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t14 92.5445
R6451 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n13 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t16 92.5445
R6452 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n14 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t49 92.5445
R6453 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n15 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t15 92.5445
R6454 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n16 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t48 92.5445
R6455 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n17 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t57 92.5445
R6456 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n18 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t58 92.5445
R6457 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n19 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t8 92.5445
R6458 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n20 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t39 92.5445
R6459 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n21 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t7 92.5445
R6460 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n23 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t17 92.5445
R6461 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n24 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t41 92.5445
R6462 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n25 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t50 92.5445
R6463 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n26 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t25 92.5445
R6464 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n28 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t29 92.5445
R6465 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n29 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t65 92.5445
R6466 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n30 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t28 92.5445
R6467 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n31 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t64 92.5445
R6468 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n32 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t10 92.5445
R6469 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n33 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t11 92.5445
R6470 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n34 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t44 92.5445
R6471 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n35 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t0 87.55
R6472 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n35 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t1 86.7044
R6473 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n35 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n49 86.4439
R6474 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n5 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n6 84.8982
R6475 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n9 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n8 84.8982
R6476 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n10 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n11 84.8982
R6477 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n14 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n13 84.8982
R6478 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n15 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n16 84.8982
R6479 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n18 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n17 84.8982
R6480 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n20 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n21 84.8982
R6481 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n24 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n23 84.8982
R6482 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n25 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n26 84.8982
R6483 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n29 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n28 84.8982
R6484 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n30 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n31 84.8982
R6485 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n33 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n32 84.8982
R6486 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n43 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t18 67.9625
R6487 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n50 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t59 67.9625
R6488 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n45 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t6 67.7525
R6489 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n52 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t45 67.7525
R6490 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n46 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n44 61.8937
R6491 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n53 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n51 61.8937
R6492 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n2 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n45 57.5119
R6493 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n3 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n43 57.5119
R6494 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n34 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n52 57.5119
R6495 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n19 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n50 57.5119
R6496 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n2 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t56 46.7545
R6497 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n3 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t21 46.7545
R6498 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n5 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t51 46.7545
R6499 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n6 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t20 46.7545
R6500 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n8 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t27 46.7545
R6501 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n9 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t63 46.7545
R6502 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n10 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t67 46.7545
R6503 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n11 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t35 46.7545
R6504 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n13 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t37 46.7545
R6505 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n14 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t13 46.7545
R6506 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n15 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t43 46.7545
R6507 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n16 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t12 46.7545
R6508 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n17 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t23 46.7545
R6509 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n18 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t24 46.7545
R6510 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n19 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t62 46.7545
R6511 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n20 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t34 46.7545
R6512 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n21 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t61 46.7545
R6513 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n23 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t9 46.7545
R6514 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n24 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t40 46.7545
R6515 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n25 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t42 46.7545
R6516 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n26 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t19 46.7545
R6517 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n28 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t22 46.7545
R6518 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n29 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t53 46.7545
R6519 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n30 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t26 46.7545
R6520 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n31 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t52 46.7545
R6521 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n32 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t66 46.7545
R6522 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n33 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t5 46.7545
R6523 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n34 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t36 46.7545
R6524 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n41 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n32 37.9969
R6525 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n40 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n30 37.9969
R6526 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n28 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n27 37.9969
R6527 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n39 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n25 37.9969
R6528 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n23 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n22 37.9969
R6529 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n20 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n42 37.9969
R6530 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n38 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n17 37.9969
R6531 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n37 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n15 37.9969
R6532 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n13 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n12 37.9969
R6533 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n36 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n10 37.9969
R6534 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n8 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n7 37.9969
R6535 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n5 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n4 37.9969
R6536 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n31 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n41 37.9654
R6537 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n40 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n29 37.9654
R6538 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n26 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n27 37.9654
R6539 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n39 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n24 37.9654
R6540 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n21 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n22 37.9654
R6541 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n42 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n19 37.9654
R6542 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n16 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n38 37.9654
R6543 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n37 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n14 37.9654
R6544 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n11 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n12 37.9654
R6545 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n36 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n9 37.9654
R6546 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n6 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n7 37.9654
R6547 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n4 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n3 37.9654
R6548 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n48 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n47 13.9641
R6549 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n55 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n54 13.9641
R6550 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n53 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n34 12.0505
R6551 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n51 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n33 12.0505
R6552 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n44 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n18 12.0505
R6553 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n46 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n2 12.0505
R6554 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n49 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t3 11.0785
R6555 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n49 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t2 11.0785
R6556 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n47 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A 9.3005
R6557 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n48 9.3005
R6558 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n54 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A 9.3005
R6559 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n55 9.3005
R6560 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n0 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n35 4.3171
R6561 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n0 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n1 3.6383
R6562 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n1 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A 3.59665
R6563 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n1 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A 3.29738
R6564 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n0 3.15388
R6565 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n0 3.03621
R6566 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n1 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A 2.99665
R6567 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n0 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A 2.97233
R6568 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n1 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A 2.688
R6569 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n0 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A 2.52972
R6570 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n0 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A 2.42304
R6571 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n1 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A 2.39665
R6572 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n0 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A 2.02323
R6573 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n1 2.01114
R6574 porb_h[0].n8 porb_h[0].n7 157.593
R6575 porb_h[0].n12 porb_h[0].n11 157.593
R6576 porb_h[0].n16 porb_h[0].n15 157.593
R6577 porb_h[0].n20 porb_h[0].n19 157.593
R6578 porb_h[0].n24 porb_h[0].n23 157.593
R6579 porb_h[0].n28 porb_h[0].n27 157.593
R6580 porb_h[0].n32 porb_h[0].n31 157.593
R6581 porb_h[0].n2 porb_h[0].n1 157.593
R6582 porb_h[0].n2 porb_h[0].n0 136.965
R6583 porb_h[0].n8 porb_h[0].n6 136.964
R6584 porb_h[0].n12 porb_h[0].n10 136.964
R6585 porb_h[0].n16 porb_h[0].n14 136.964
R6586 porb_h[0].n20 porb_h[0].n18 136.964
R6587 porb_h[0].n24 porb_h[0].n22 136.964
R6588 porb_h[0].n28 porb_h[0].n26 136.964
R6589 porb_h[0].n32 porb_h[0].n30 136.964
R6590 porb_h[0].n6 porb_h[0].t9 21.2805
R6591 porb_h[0].n6 porb_h[0].t8 21.2805
R6592 porb_h[0].n10 porb_h[0].t4 21.2805
R6593 porb_h[0].n10 porb_h[0].t14 21.2805
R6594 porb_h[0].n14 porb_h[0].t5 21.2805
R6595 porb_h[0].n14 porb_h[0].t13 21.2805
R6596 porb_h[0].n18 porb_h[0].t0 21.2805
R6597 porb_h[0].n18 porb_h[0].t6 21.2805
R6598 porb_h[0].n22 porb_h[0].t7 21.2805
R6599 porb_h[0].n22 porb_h[0].t1 21.2805
R6600 porb_h[0].n26 porb_h[0].t3 21.2805
R6601 porb_h[0].n26 porb_h[0].t11 21.2805
R6602 porb_h[0].n30 porb_h[0].t12 21.2805
R6603 porb_h[0].n30 porb_h[0].t10 21.2805
R6604 porb_h[0].n0 porb_h[0].t2 21.2805
R6605 porb_h[0].n0 porb_h[0].t15 21.2805
R6606 porb_h[0].n7 porb_h[0].t30 17.8272
R6607 porb_h[0].n7 porb_h[0].t29 17.8272
R6608 porb_h[0].n11 porb_h[0].t26 17.8272
R6609 porb_h[0].n11 porb_h[0].t25 17.8272
R6610 porb_h[0].n15 porb_h[0].t28 17.8272
R6611 porb_h[0].n15 porb_h[0].t24 17.8272
R6612 porb_h[0].n19 porb_h[0].t19 17.8272
R6613 porb_h[0].n19 porb_h[0].t27 17.8272
R6614 porb_h[0].n23 porb_h[0].t22 17.8272
R6615 porb_h[0].n23 porb_h[0].t17 17.8272
R6616 porb_h[0].n27 porb_h[0].t18 17.8272
R6617 porb_h[0].n27 porb_h[0].t23 17.8272
R6618 porb_h[0].n31 porb_h[0].t16 17.8272
R6619 porb_h[0].n31 porb_h[0].t31 17.8272
R6620 porb_h[0].n1 porb_h[0].t21 17.8272
R6621 porb_h[0].n1 porb_h[0].t20 17.8272
R6622 porb_h[0].n9 porb_h[0].n8 9.98018
R6623 porb_h[0].n13 porb_h[0].n12 9.98018
R6624 porb_h[0].n17 porb_h[0].n16 9.98018
R6625 porb_h[0].n21 porb_h[0].n20 9.98018
R6626 porb_h[0].n25 porb_h[0].n24 9.98018
R6627 porb_h[0].n29 porb_h[0].n28 9.98018
R6628 porb_h[0].n33 porb_h[0].n32 9.98018
R6629 porb_h[0].n3 porb_h[0].n2 9.98018
R6630 porb_h[0] porb_h[0].n33 2.80521
R6631 porb_h[0].n33 porb_h[0].n29 0.402562
R6632 porb_h[0].n29 porb_h[0].n25 0.402562
R6633 porb_h[0].n25 porb_h[0].n21 0.402562
R6634 porb_h[0].n21 porb_h[0].n17 0.402562
R6635 porb_h[0].n17 porb_h[0].n13 0.402562
R6636 porb_h[0].n13 porb_h[0].n9 0.402562
R6637 porb_h[0].n9 porb_h[0].n5 0.314933
R6638 porb_h[0].n4 porb_h[0] 0.213735
R6639 porb_h[0].n5 porb_h[0].n4 0.143882
R6640 porb_h[0].n5 porb_h[0] 0.1255
R6641 porb_h[0].n4 porb_h[0].n3 0.0793043
R6642 porb_h[0].n3 porb_h[0] 0.0793043
R6643 avdd.n450 avdd.n449 85267.4
R6644 avdd.n451 avdd.n450 81309.1
R6645 avdd.n451 avdd.n118 80879.3
R6646 avdd.n448 avdd.n117 73784.8
R6647 avdd.n122 avdd.n118 72120.8
R6648 avdd.n452 avdd.n117 70431.9
R6649 avdd.n452 avdd.n116 54951.4
R6650 avdd.n123 avdd.n116 46015.8
R6651 avdd.n121 avdd.n119 34238.3
R6652 avdd.n448 avdd.n120 31085.1
R6653 avdd.n122 avdd.n121 29064.7
R6654 avdd.n123 avdd.n120 18756.4
R6655 avdd.n449 avdd.n119 3423.96
R6656 avdd.n431 avdd.n396 2710.45
R6657 avdd.n431 avdd.n397 2710.45
R6658 avdd.n446 avdd.n114 2105.51
R6659 avdd.n455 avdd.n454 1951.99
R6660 avdd.n490 avdd.n486 1643.17
R6661 avdd.n524 avdd.n466 1643.17
R6662 avdd.n524 avdd.n467 1643.17
R6663 avdd.n513 avdd.n477 1643.17
R6664 avdd.n504 avdd.n477 1643.17
R6665 avdd.n521 avdd.n468 1643.17
R6666 avdd.n102 avdd.n97 1544.9
R6667 avdd.n90 avdd.n44 1544.9
R6668 avdd.n91 avdd.n44 1544.9
R6669 avdd.n195 avdd.n186 1483.97
R6670 avdd.n192 avdd.n186 1483.97
R6671 avdd.n205 avdd.n179 1483.97
R6672 avdd.n203 avdd.n179 1483.97
R6673 avdd.n154 avdd.n146 1405.34
R6674 avdd.n150 avdd.n146 1405.34
R6675 avdd.n168 avdd.n136 1405.34
R6676 avdd.n168 avdd.n137 1405.34
R6677 avdd.n453 avdd.n115 1333.59
R6678 avdd.n421 avdd.n397 1322.79
R6679 avdd.n82 avdd.n50 1250.07
R6680 avdd.n83 avdd.n50 1250.07
R6681 avdd.n83 avdd.n49 1250.07
R6682 avdd.n82 avdd.n49 1250.07
R6683 avdd.n405 avdd.n396 1232.38
R6684 avdd.n415 avdd.n406 1210.76
R6685 avdd.n424 avdd.n422 1210.76
R6686 avdd.n15 avdd.n14 1151.79
R6687 avdd.n29 avdd.n4 1151.79
R6688 avdd.n441 avdd.n440 1132.55
R6689 avdd.n46 avdd.n42 1126.24
R6690 avdd.n47 avdd.n46 1126.24
R6691 avdd.n104 avdd.n38 1126.24
R6692 avdd.n104 avdd.n39 1126.24
R6693 avdd.n73 avdd.n57 1110.52
R6694 avdd.n73 avdd.n58 1110.52
R6695 avdd.n76 avdd.n57 1110.52
R6696 avdd.n76 avdd.n58 1110.52
R6697 avdd.n490 avdd.n482 1106.59
R6698 avdd.n482 avdd.n466 1106.59
R6699 avdd.n484 avdd.n483 1106.59
R6700 avdd.n483 avdd.n467 1106.59
R6701 avdd.n502 avdd.n501 1106.59
R6702 avdd.n501 avdd.n476 1106.59
R6703 avdd.n520 avdd.n519 1106.59
R6704 avdd.n519 avdd.n470 1106.59
R6705 avdd.n405 avdd.n404 955.241
R6706 avdd.n421 avdd.n399 955.241
R6707 avdd.n196 avdd.n185 910.034
R6708 avdd.n185 avdd.n182 910.034
R6709 avdd.n183 avdd.n178 910.034
R6710 avdd.n183 avdd.n180 910.034
R6711 avdd.n151 avdd.n143 831.414
R6712 avdd.n151 avdd.n142 831.414
R6713 avdd.n165 avdd.n138 831.414
R6714 avdd.n165 avdd.n139 831.414
R6715 avdd.n447 avdd.n445 806.308
R6716 avdd.n404 avdd.n403 733.139
R6717 avdd.n416 avdd.n403 733.139
R6718 avdd.n406 avdd.n405 733.139
R6719 avdd.n428 avdd.n399 733.139
R6720 avdd.n428 avdd.n400 733.139
R6721 avdd.n422 avdd.n421 733.139
R6722 avdd.n21 avdd.n11 733.139
R6723 avdd.n11 avdd.n9 733.139
R6724 avdd.n6 avdd.n3 733.139
R6725 avdd.n7 avdd.n6 733.139
R6726 avdd.n491 avdd.t118 673.615
R6727 avdd.n491 avdd.t116 673.615
R6728 avdd.n523 avdd.t116 673.615
R6729 avdd.n522 avdd.t20 673.615
R6730 avdd.n196 avdd.n195 573.932
R6731 avdd.n197 avdd.n196 573.932
R6732 avdd.n197 avdd.n178 573.932
R6733 avdd.n205 avdd.n178 573.932
R6734 avdd.n192 avdd.n182 573.932
R6735 avdd.n199 avdd.n182 573.932
R6736 avdd.n199 avdd.n180 573.932
R6737 avdd.n203 avdd.n180 573.932
R6738 avdd.n154 avdd.n143 573.932
R6739 avdd.n159 avdd.n143 573.932
R6740 avdd.n159 avdd.n138 573.932
R6741 avdd.n138 avdd.n136 573.932
R6742 avdd.n150 avdd.n142 573.932
R6743 avdd.n161 avdd.n142 573.932
R6744 avdd.n161 avdd.n139 573.932
R6745 avdd.n139 avdd.n137 573.932
R6746 avdd.n492 avdd.n482 536.587
R6747 avdd.n492 avdd.n483 536.587
R6748 avdd.n513 avdd.n476 536.587
R6749 avdd.n520 avdd.n469 536.587
R6750 avdd.n502 avdd.n469 536.587
R6751 avdd.n504 avdd.n502 536.587
R6752 avdd.n473 avdd.n470 536.587
R6753 avdd.n515 avdd.n470 536.587
R6754 avdd.n515 avdd.n476 536.587
R6755 avdd.n521 avdd.n520 536.587
R6756 avdd.n404 avdd.n398 522.828
R6757 avdd.n486 avdd.n485 488.151
R6758 avdd.n473 avdd.n472 488.151
R6759 avdd.n416 avdd.n415 477.622
R6760 avdd.n417 avdd.n416 477.622
R6761 avdd.n417 avdd.n400 477.622
R6762 avdd.n424 avdd.n400 477.622
R6763 avdd.n444 avdd.n124 446.837
R6764 avdd.n503 avdd.t20 442.757
R6765 avdd.n514 avdd.t20 442.757
R6766 avdd.n399 avdd.n398 432.414
R6767 avdd.n90 avdd.n47 418.656
R6768 avdd.n47 avdd.n41 418.656
R6769 avdd.n41 avdd.n39 418.656
R6770 avdd.n98 avdd.n39 418.656
R6771 avdd.n91 avdd.n42 418.656
R6772 avdd.n95 avdd.n42 418.656
R6773 avdd.n95 avdd.n38 418.656
R6774 avdd.n102 avdd.n38 418.656
R6775 avdd.n21 avdd.n20 418.656
R6776 avdd.n22 avdd.n21 418.656
R6777 avdd.n22 avdd.n3 418.656
R6778 avdd.n29 avdd.n3 418.656
R6779 avdd.n14 avdd.n9 418.656
R6780 avdd.n23 avdd.n9 418.656
R6781 avdd.n23 avdd.n7 418.656
R6782 avdd.n27 avdd.n7 418.656
R6783 avdd.n523 avdd.n522 335.014
R6784 avdd.n285 avdd.n277 321.882
R6785 avdd.n290 avdd.n277 321.882
R6786 avdd.n290 avdd.n270 321.882
R6787 avdd.n301 avdd.n270 321.882
R6788 avdd.n302 avdd.n301 321.882
R6789 avdd.n302 avdd.n268 321.882
R6790 avdd.n307 avdd.n268 321.882
R6791 avdd.n307 avdd.n259 321.882
R6792 avdd.n324 avdd.n259 321.882
R6793 avdd.n324 avdd.n258 321.882
R6794 avdd.n329 avdd.n258 321.882
R6795 avdd.n329 avdd.n239 321.882
R6796 avdd.n338 avdd.n239 321.882
R6797 avdd.n338 avdd.n237 321.882
R6798 avdd.n342 avdd.n237 321.882
R6799 avdd.n343 avdd.n342 321.882
R6800 avdd.n343 avdd.n217 321.882
R6801 avdd.n218 avdd.n217 321.882
R6802 avdd.n219 avdd.n218 321.882
R6803 avdd.n348 avdd.n219 321.882
R6804 avdd.n348 avdd.n227 321.882
R6805 avdd.n228 avdd.n227 321.882
R6806 avdd.n352 avdd.n228 321.882
R6807 avdd.n352 avdd.n235 321.882
R6808 avdd.n236 avdd.n235 321.882
R6809 avdd.n356 avdd.n236 321.882
R6810 avdd.n147 avdd.n119 303.062
R6811 avdd.n286 avdd.n278 301.973
R6812 avdd.n202 avdd.n177 288.753
R6813 avdd.n191 avdd.n190 288.753
R6814 avdd.t11 avdd.n73 281.277
R6815 avdd.n356 avdd.t48 280.652
R6816 avdd.n498 avdd.n497 277.113
R6817 avdd.n359 avdd.t49 275.541
R6818 avdd.n358 avdd.t58 275.539
R6819 avdd.n280 avdd.t35 274.385
R6820 avdd.n281 avdd.t50 274.384
R6821 avdd.n419 avdd.n395 257.882
R6822 avdd.n487 avdd.n478 255.095
R6823 avdd.n75 avdd.t23 254.85
R6824 avdd.t26 avdd.n51 251.358
R6825 avdd.t26 avdd.n52 251.358
R6826 avdd.n410 avdd.n394 240.565
R6827 avdd.n425 avdd.n420 236.424
R6828 avdd.n412 avdd.n411 236.424
R6829 avdd.t28 avdd.n397 227.356
R6830 avdd.n26 avdd.n2 225.13
R6831 avdd.n16 avdd.n13 225.13
R6832 avdd.n493 avdd.t119 222.696
R6833 avdd.n474 avdd.t110 222.696
R6834 avdd.n527 avdd.t117 222.696
R6835 avdd.n54 avdd.t24 222.696
R6836 avdd.n69 avdd.t12 222.696
R6837 avdd.t6 avdd.n396 214.845
R6838 avdd.n494 avdd.n478 211.953
R6839 avdd.n495 avdd.n494 211.953
R6840 avdd.n432 avdd.n395 211.298
R6841 avdd.n433 avdd.n394 205.964
R6842 avdd.n518 avdd.n471 205.554
R6843 avdd.n518 avdd.n517 205.554
R6844 avdd.n500 avdd.n499 205.554
R6845 avdd.n500 avdd.n475 205.554
R6846 avdd.n496 avdd.n495 205.554
R6847 avdd.t14 avdd.n10 203.571
R6848 avdd.t8 avdd.n10 203.571
R6849 avdd.t8 avdd.n5 203.571
R6850 avdd.t13 avdd.n5 203.571
R6851 avdd.n168 avdd.t114 201.782
R6852 avdd.n106 avdd.t124 192.494
R6853 avdd.n206 avdd.n177 191.774
R6854 avdd.n190 avdd.n189 191.774
R6855 avdd.n106 avdd.t123 191.234
R6856 avdd.t80 avdd.n186 187.776
R6857 avdd.t90 avdd.n179 187.776
R6858 avdd.n285 avdd.n284 185
R6859 avdd.n277 avdd.n276 185
R6860 avdd.n287 avdd.n277 185
R6861 avdd.n291 avdd.n290 185
R6862 avdd.n290 avdd.n289 185
R6863 avdd.n271 avdd.n270 185
R6864 avdd.n288 avdd.n270 185
R6865 avdd.n301 avdd.n300 185
R6866 avdd.n301 avdd.n269 185
R6867 avdd.n302 avdd.n267 185
R6868 avdd.n303 avdd.n302 185
R6869 avdd.n309 avdd.n268 185
R6870 avdd.n304 avdd.n268 185
R6871 avdd.n308 avdd.n307 185
R6872 avdd.n307 avdd.n306 185
R6873 avdd.n260 avdd.n259 185
R6874 avdd.n305 avdd.n259 185
R6875 avdd.n324 avdd.n323 185
R6876 avdd.n325 avdd.n324 185
R6877 avdd.n258 avdd.n257 185
R6878 avdd.n326 avdd.n258 185
R6879 avdd.n330 avdd.n329 185
R6880 avdd.n329 avdd.n328 185
R6881 avdd.n240 avdd.n239 185
R6882 avdd.n327 avdd.n239 185
R6883 avdd.n338 avdd.n337 185
R6884 avdd.n339 avdd.n338 185
R6885 avdd.n241 avdd.n237 185
R6886 avdd.n340 avdd.n237 185
R6887 avdd.n342 avdd.n238 185
R6888 avdd.n342 avdd.n341 185
R6889 avdd.n343 avdd.n216 185
R6890 avdd.n344 avdd.n343 185
R6891 avdd.n379 avdd.n217 185
R6892 avdd.n345 avdd.n217 185
R6893 avdd.n378 avdd.n218 185
R6894 avdd.n346 avdd.n218 185
R6895 avdd.n377 avdd.n219 185
R6896 avdd.n347 avdd.n219 185
R6897 avdd.n348 avdd.n220 185
R6898 avdd.n349 avdd.n348 185
R6899 avdd.n371 avdd.n227 185
R6900 avdd.n350 avdd.n227 185
R6901 avdd.n370 avdd.n228 185
R6902 avdd.n351 avdd.n228 185
R6903 avdd.n352 avdd.n229 185
R6904 avdd.n353 avdd.n352 185
R6905 avdd.n364 avdd.n235 185
R6906 avdd.n354 avdd.n235 185
R6907 avdd.n363 avdd.n236 185
R6908 avdd.n355 avdd.n236 185
R6909 avdd.n362 avdd.n356 185
R6910 avdd.t102 avdd.n147 184.964
R6911 avdd.t104 avdd.n152 184.964
R6912 avdd.n152 avdd.t108 184.964
R6913 avdd.n166 avdd.t106 184.964
R6914 avdd.t78 avdd.n166 184.964
R6915 avdd.n410 avdd.n409 182.965
R6916 avdd.n419 avdd.n401 182.965
R6917 avdd.n15 avdd.n12 180.113
R6918 avdd.n28 avdd.n4 180.113
R6919 avdd.n201 avdd.n176 178.825
R6920 avdd.n187 avdd.n181 178.825
R6921 avdd.n207 avdd.n176 172.8
R6922 avdd.n188 avdd.n187 172.8
R6923 avdd.t21 avdd.n193 172.359
R6924 avdd.n193 avdd.t0 172.359
R6925 avdd.t2 avdd.n184 172.359
R6926 avdd.n184 avdd.t88 172.359
R6927 avdd.n144 avdd.n141 163.766
R6928 avdd.n164 avdd.n163 163.766
R6929 avdd.n30 avdd.n2 159.016
R6930 avdd.n19 avdd.n16 159.016
R6931 avdd.n156 avdd.n144 158.494
R6932 avdd.n164 avdd.n140 158.494
R6933 avdd.n169 avdd.n135 156.606
R6934 avdd.n52 avdd.n45 154.582
R6935 avdd.n100 avdd.n99 154.055
R6936 avdd.n367 avdd.n233 151.065
R6937 avdd.n374 avdd.n225 151.065
R6938 avdd.n251 avdd.n248 151.065
R6939 avdd.n334 avdd.n255 151.065
R6940 avdd.n320 avdd.n319 151.065
R6941 avdd.n312 avdd.n264 151.065
R6942 avdd.n297 avdd.n273 151.065
R6943 avdd.n231 avdd.n230 151.065
R6944 avdd.n223 avdd.n222 151.065
R6945 avdd.n246 avdd.n245 151.065
R6946 avdd.n244 avdd.n243 151.065
R6947 avdd.n317 avdd.n316 151.065
R6948 avdd.n263 avdd.n262 151.065
R6949 avdd.n294 avdd.n293 151.065
R6950 avdd.n149 avdd.n148 149.828
R6951 avdd.t94 avdd.n45 145.159
R6952 avdd.t94 avdd.n40 145.159
R6953 avdd.t9 avdd.n40 145.159
R6954 avdd.n103 avdd.t9 145.159
R6955 avdd.n103 avdd.t111 145.159
R6956 avdd.n427 avdd.n401 144.941
R6957 avdd.n427 avdd.n426 144.941
R6958 avdd.n409 avdd.n407 144.941
R6959 avdd.n407 avdd.n402 144.941
R6960 avdd.n420 avdd.n419 144.941
R6961 avdd.n411 avdd.n410 144.941
R6962 avdd.n25 avdd.n1 144.941
R6963 avdd.n17 avdd.n8 144.941
R6964 avdd.n31 avdd.n1 143.435
R6965 avdd.n18 avdd.n17 143.435
R6966 avdd.t34 avdd.n286 141.143
R6967 avdd.n97 avdd.n96 139.143
R6968 avdd.t18 avdd.n62 122.499
R6969 avdd.n63 avdd.t18 122.436
R6970 avdd.n75 avdd.n51 121.903
R6971 avdd.n71 avdd.n70 120.526
R6972 avdd.n393 avdd.t93 116.66
R6973 avdd.n387 avdd.t29 116.1
R6974 avdd.n392 avdd.t7 115.799
R6975 avdd avdd.t15 113.477
R6976 avdd.n89 avdd.n86 111.49
R6977 avdd.n65 avdd.t27 111.349
R6978 avdd.n84 avdd.n48 110.823
R6979 avdd.n191 avdd.n181 109.93
R6980 avdd.n200 avdd.n181 109.93
R6981 avdd.n201 avdd.n200 109.93
R6982 avdd.n202 avdd.n201 109.93
R6983 avdd.n149 avdd.n141 109.93
R6984 avdd.n162 avdd.n141 109.93
R6985 avdd.n163 avdd.n162 109.93
R6986 avdd.n163 avdd.n135 109.93
R6987 avdd.t82 avdd.n413 109.373
R6988 avdd.n289 avdd.n287 104.349
R6989 avdd.n303 avdd.n269 104.349
R6990 avdd.n306 avdd.n304 104.349
R6991 avdd.n326 avdd.n325 104.349
R6992 avdd.n328 avdd.n327 104.349
R6993 avdd.n341 avdd.n340 104.349
R6994 avdd.n346 avdd.n345 104.349
R6995 avdd.n349 avdd.n347 104.349
R6996 avdd.n353 avdd.n351 104.349
R6997 avdd.n355 avdd.n354 104.349
R6998 avdd.n70 avdd.n48 103.529
R6999 avdd.n512 avdd.n511 103.234
R7000 avdd.n86 avdd.n84 103.233
R7001 avdd.n389 avdd.n388 101.951
R7002 avdd.n391 avdd.n390 101.942
R7003 avdd.n387 avdd.n386 101.936
R7004 avdd.n409 avdd.n408 100.141
R7005 avdd.n288 avdd.t55 100.001
R7006 avdd.t64 avdd.n344 100.001
R7007 avdd.n105 avdd.n37 99.8235
R7008 avdd.n88 avdd.n35 99.2229
R7009 avdd.n128 avdd.t103 97.5645
R7010 avdd.n128 avdd.t105 97.4016
R7011 avdd.n131 avdd.t79 97.3968
R7012 avdd.n132 avdd.t115 97.392
R7013 avdd.n129 avdd.t109 97.392
R7014 avdd.n130 avdd.t107 97.3758
R7015 avdd.t92 avdd.t86 96.1629
R7016 avdd.n339 avdd.t66 95.6527
R7017 avdd.n74 avdd.t11 94.5219
R7018 avdd.t23 avdd.n74 94.5219
R7019 avdd.n412 avdd.n402 91.4829
R7020 avdd.n418 avdd.n402 91.4829
R7021 avdd.n426 avdd.n418 91.4829
R7022 avdd.n426 avdd.n425 91.4829
R7023 avdd.n510 avdd.n505 89.9697
R7024 avdd.n305 avdd.t53 86.957
R7025 avdd.t36 avdd.n350 86.957
R7026 avdd.n101 avdd.n100 85.9071
R7027 avdd.t84 avdd.n423 85.0672
R7028 avdd.n61 avdd.t17 82.9645
R7029 avdd.n414 avdd.t4 82.9538
R7030 avdd.n60 avdd.t19 82.8472
R7031 avdd.n408 avdd.n401 82.824
R7032 avdd.n494 avdd.n493 82.6717
R7033 avdd.t68 avdd.n305 82.6092
R7034 avdd.n350 avdd.t38 82.6092
R7035 avdd.n170 avdd.n134 82.4166
R7036 avdd.n155 avdd.n145 81.4941
R7037 avdd.n89 avdd.n88 80.1887
R7038 avdd.n88 avdd.n87 80.1887
R7039 avdd.n87 avdd.n37 80.1887
R7040 avdd.n99 avdd.n37 80.1887
R7041 avdd.n13 avdd.n8 80.1887
R7042 avdd.n24 avdd.n8 80.1887
R7043 avdd.n25 avdd.n24 80.1887
R7044 avdd.n26 avdd.n25 80.1887
R7045 avdd.n517 avdd.n474 77.3594
R7046 avdd.n210 avdd.n125 75.8935
R7047 avdd.n174 avdd.n126 75.8557
R7048 avdd.n173 avdd.n127 75.8402
R7049 avdd.n286 avdd.n285 74.7887
R7050 avdd.t62 avdd.n339 73.9135
R7051 avdd.t96 avdd.t97 71.8581
R7052 avdd.n497 avdd.n496 70.5901
R7053 avdd.n71 avdd.n69 70.3317
R7054 avdd.t40 avdd.n288 69.5657
R7055 avdd.n344 avdd.t30 69.5657
R7056 avdd.n153 avdd.t102 68.602
R7057 avdd.n153 avdd.t104 68.602
R7058 avdd.n160 avdd.t108 68.602
R7059 avdd.n160 avdd.t106 68.602
R7060 avdd.n167 avdd.t78 68.602
R7061 avdd.t114 avdd.n167 68.602
R7062 avdd.n489 avdd.n487 65.8738
R7063 avdd.n194 avdd.t80 63.9272
R7064 avdd.n194 avdd.t21 63.9272
R7065 avdd.n198 avdd.t0 63.9272
R7066 avdd.n198 avdd.t2 63.9272
R7067 avdd.n204 avdd.t88 63.9272
R7068 avdd.n204 avdd.t90 63.9272
R7069 avdd.n61 avdd.t16 61.2493
R7070 avdd.n527 avdd.n526 61.1697
R7071 avdd.t42 avdd.n303 60.8701
R7072 avdd.t32 avdd.n346 60.8701
R7073 avdd.n56 avdd.n54 60.1321
R7074 avdd.n34 avdd.t95 60.1061
R7075 avdd.n35 avdd.t10 60.1061
R7076 avdd.n105 avdd.t112 60.1061
R7077 avdd.t100 avdd.n429 58.649
R7078 avdd.n430 avdd.t100 57.5923
R7079 avdd.n429 avdd.t97 56.5355
R7080 avdd.n328 avdd.t44 56.5222
R7081 avdd.n354 avdd.t51 56.5222
R7082 avdd.t44 avdd.n326 47.8266
R7083 avdd.t51 avdd.n353 47.8266
R7084 avdd.n102 avdd.n101 46.2505
R7085 avdd.t111 avdd.n102 46.2505
R7086 avdd.n95 avdd.n94 46.2505
R7087 avdd.t9 avdd.n95 46.2505
R7088 avdd.n92 avdd.n91 46.2505
R7089 avdd.n91 avdd.t94 46.2505
R7090 avdd.n99 avdd.n98 46.2505
R7091 avdd.n87 avdd.n41 46.2505
R7092 avdd.t9 avdd.n41 46.2505
R7093 avdd.n90 avdd.n89 46.2505
R7094 avdd.t94 avdd.n90 46.2505
R7095 avdd.n27 avdd.n26 46.2505
R7096 avdd.n24 avdd.n23 46.2505
R7097 avdd.n23 avdd.t8 46.2505
R7098 avdd.n14 avdd.n13 46.2505
R7099 avdd.n14 avdd.t14 46.2505
R7100 avdd.n30 avdd.n29 46.2505
R7101 avdd.n29 avdd.t13 46.2505
R7102 avdd.n22 avdd.n0 46.2505
R7103 avdd.t8 avdd.n22 46.2505
R7104 avdd.n20 avdd.n19 46.2505
R7105 avdd.t4 avdd.t113 45.4399
R7106 avdd.n93 avdd.n35 45.2587
R7107 avdd.n105 avdd.n36 45.1595
R7108 avdd.n304 avdd.t42 43.4788
R7109 avdd.n347 avdd.t32 43.4788
R7110 avdd.n517 avdd.n516 43.4342
R7111 avdd.n516 avdd.n475 43.4342
R7112 avdd.n512 avdd.n475 43.4342
R7113 avdd.t96 avdd.t84 43.3264
R7114 avdd.n98 avdd.n96 40.8622
R7115 avdd.n20 avdd.n12 37.5124
R7116 avdd.n28 avdd.n27 37.5124
R7117 avdd.n82 avdd.n81 37.0005
R7118 avdd.t26 avdd.n82 37.0005
R7119 avdd.n84 avdd.n83 37.0005
R7120 avdd.n83 avdd.t26 37.0005
R7121 avdd.n425 avdd.n424 37.0005
R7122 avdd.n424 avdd.t96 37.0005
R7123 avdd.n418 avdd.n417 37.0005
R7124 avdd.n417 avdd.t113 37.0005
R7125 avdd.n415 avdd.n412 37.0005
R7126 avdd.n415 avdd.t92 37.0005
R7127 avdd.n284 avdd.n278 36.1417
R7128 avdd.n284 avdd.n276 36.1417
R7129 avdd.n291 avdd.n276 36.1417
R7130 avdd.n291 avdd.n271 36.1417
R7131 avdd.n300 avdd.n271 36.1417
R7132 avdd.n300 avdd.n267 36.1417
R7133 avdd.n309 avdd.n267 36.1417
R7134 avdd.n309 avdd.n308 36.1417
R7135 avdd.n308 avdd.n260 36.1417
R7136 avdd.n323 avdd.n260 36.1417
R7137 avdd.n323 avdd.n257 36.1417
R7138 avdd.n330 avdd.n257 36.1417
R7139 avdd.n330 avdd.n240 36.1417
R7140 avdd.n337 avdd.n240 36.1417
R7141 avdd.n337 avdd.n241 36.1417
R7142 avdd.n241 avdd.n238 36.1417
R7143 avdd.n238 avdd.n216 36.1417
R7144 avdd.n379 avdd.n216 36.1417
R7145 avdd.n379 avdd.n378 36.1417
R7146 avdd.n378 avdd.n377 36.1417
R7147 avdd.n377 avdd.n220 36.1417
R7148 avdd.n371 avdd.n220 36.1417
R7149 avdd.n371 avdd.n370 36.1417
R7150 avdd.n370 avdd.n229 36.1417
R7151 avdd.n364 avdd.n229 36.1417
R7152 avdd.n364 avdd.n363 36.1417
R7153 avdd.n363 avdd.n362 36.1417
R7154 avdd.n289 avdd.t40 34.7831
R7155 avdd.n341 avdd.t30 34.7831
R7156 avdd.n456 avdd.n113 32.8461
R7157 avdd.t86 avdd.n414 32.2308
R7158 avdd.n499 avdd.n498 32.2138
R7159 avdd.n505 avdd.n499 32.2138
R7160 avdd.n70 avdd.n58 30.8338
R7161 avdd.n74 avdd.n58 30.8338
R7162 avdd.n57 avdd.n53 30.8338
R7163 avdd.n74 avdd.n57 30.8338
R7164 avdd.n203 avdd.n202 30.8338
R7165 avdd.n204 avdd.n203 30.8338
R7166 avdd.n200 avdd.n199 30.8338
R7167 avdd.n199 avdd.n198 30.8338
R7168 avdd.n192 avdd.n191 30.8338
R7169 avdd.n194 avdd.n192 30.8338
R7170 avdd.n206 avdd.n205 30.8338
R7171 avdd.n205 avdd.n204 30.8338
R7172 avdd.n197 avdd.n175 30.8338
R7173 avdd.n198 avdd.n197 30.8338
R7174 avdd.n195 avdd.n189 30.8338
R7175 avdd.n195 avdd.n194 30.8338
R7176 avdd.n137 avdd.n135 30.8338
R7177 avdd.n167 avdd.n137 30.8338
R7178 avdd.n162 avdd.n161 30.8338
R7179 avdd.n161 avdd.n160 30.8338
R7180 avdd.n150 avdd.n149 30.8338
R7181 avdd.n153 avdd.n150 30.8338
R7182 avdd.n136 avdd.n134 30.8338
R7183 avdd.n167 avdd.n136 30.8338
R7184 avdd.n159 avdd.n158 30.8338
R7185 avdd.n160 avdd.n159 30.8338
R7186 avdd.n155 avdd.n154 30.8338
R7187 avdd.n154 avdd.n153 30.8338
R7188 avdd.n156 avdd.n155 30.6366
R7189 avdd.n158 avdd.n156 30.6366
R7190 avdd.n140 avdd.n134 30.6366
R7191 avdd.n287 avdd.t34 30.4353
R7192 avdd.n340 avdd.t62 30.4353
R7193 avdd.n531 avdd.n461 30.3507
R7194 avdd.n423 avdd.t28 30.1173
R7195 avdd.n487 avdd.n486 29.9905
R7196 avdd.n157 avdd.n140 29.7972
R7197 avdd.n526 avdd.n465 27.7338
R7198 avdd.n59 avdd.n53 26.5298
R7199 avdd.n532 avdd.n531 26.4883
R7200 avdd.n474 avdd.n473 26.4291
R7201 avdd.n516 avdd.n515 26.4291
R7202 avdd.n515 avdd.n514 26.4291
R7203 avdd.n513 avdd.n512 26.4291
R7204 avdd.n514 avdd.n513 26.4291
R7205 avdd.n498 avdd.n469 26.4291
R7206 avdd.n503 avdd.n469 26.4291
R7207 avdd.n505 avdd.n504 26.4291
R7208 avdd.n504 avdd.n503 26.4291
R7209 avdd.n521 avdd.n462 26.4291
R7210 avdd.n522 avdd.n521 26.4291
R7211 avdd.n525 avdd.n524 26.4291
R7212 avdd.n524 avdd.n523 26.4291
R7213 avdd.n493 avdd.n492 26.4291
R7214 avdd.n492 avdd.n491 26.4291
R7215 avdd.n73 avdd.n72 26.4291
R7216 avdd.n77 avdd.n76 26.4291
R7217 avdd.n76 avdd.n75 26.4291
R7218 avdd.n506 avdd.n461 24.7038
R7219 avdd.n488 avdd.n460 23.9714
R7220 avdd.n457 avdd.n456 23.8601
R7221 avdd.n496 avdd.n465 23.4672
R7222 avdd.n306 avdd.t68 21.7396
R7223 avdd.t38 avdd.n349 21.7396
R7224 avdd.n489 avdd.n488 19.7047
R7225 avdd.t92 avdd.t82 19.0216
R7226 avdd.n189 avdd.n188 18.9731
R7227 avdd.n188 avdd.n175 18.9731
R7228 avdd.n207 avdd.n206 18.9731
R7229 avdd.n55 avdd.n49 18.5005
R7230 avdd.n51 avdd.n49 18.5005
R7231 avdd.n64 avdd.n50 18.5005
R7232 avdd.n52 avdd.n50 18.5005
R7233 avdd.n397 avdd.n395 18.5005
R7234 avdd.n407 avdd.n403 18.5005
R7235 avdd.n414 avdd.n403 18.5005
R7236 avdd.n428 avdd.n427 18.5005
R7237 avdd.n429 avdd.n428 18.5005
R7238 avdd.n422 avdd.n420 18.5005
R7239 avdd.n423 avdd.n422 18.5005
R7240 avdd.n411 avdd.n406 18.5005
R7241 avdd.n413 avdd.n406 18.5005
R7242 avdd.n396 avdd.n394 18.5005
R7243 avdd.n17 avdd.n11 18.5005
R7244 avdd.n11 avdd.n10 18.5005
R7245 avdd.n6 avdd.n1 18.5005
R7246 avdd.n6 avdd.n5 18.5005
R7247 avdd.n4 avdd.n2 18.5005
R7248 avdd.n16 avdd.n15 18.5005
R7249 avdd.n208 avdd.n207 18.1934
R7250 avdd.n488 avdd.n481 18.0934
R7251 avdd.n233 avdd.t74 17.8272
R7252 avdd.n233 avdd.t52 17.8272
R7253 avdd.n225 avdd.t33 17.8272
R7254 avdd.n225 avdd.t70 17.8272
R7255 avdd.n248 avdd.t31 17.8272
R7256 avdd.n248 avdd.t65 17.8272
R7257 avdd.n255 avdd.t67 17.8272
R7258 avdd.n255 avdd.t63 17.8272
R7259 avdd.n319 avdd.t54 17.8272
R7260 avdd.n319 avdd.t45 17.8272
R7261 avdd.n264 avdd.t76 17.8272
R7262 avdd.n264 avdd.t69 17.8272
R7263 avdd.n273 avdd.t75 17.8272
R7264 avdd.n273 avdd.t56 17.8272
R7265 avdd.n230 avdd.t37 17.8272
R7266 avdd.n230 avdd.t59 17.8272
R7267 avdd.n222 avdd.t47 17.8272
R7268 avdd.n222 avdd.t39 17.8272
R7269 avdd.n245 avdd.t46 17.8272
R7270 avdd.n245 avdd.t72 17.8272
R7271 avdd.n243 avdd.t73 17.8272
R7272 avdd.n243 avdd.t71 17.8272
R7273 avdd.n316 avdd.t60 17.8272
R7274 avdd.n316 avdd.t57 17.8272
R7275 avdd.n262 avdd.t43 17.8272
R7276 avdd.n262 avdd.t77 17.8272
R7277 avdd.n293 avdd.t41 17.8272
R7278 avdd.n293 avdd.t61 17.8272
R7279 avdd.n325 avdd.t53 17.3918
R7280 avdd.n351 avdd.t36 17.3918
R7281 avdd.n55 avdd.n48 17.1773
R7282 avdd.n151 avdd.n144 16.8187
R7283 avdd.n152 avdd.n151 16.8187
R7284 avdd.n165 avdd.n164 16.8187
R7285 avdd.n166 avdd.n165 16.8187
R7286 avdd.n148 avdd.n146 16.8187
R7287 avdd.n147 avdd.n146 16.8187
R7288 avdd.n169 avdd.n168 16.8187
R7289 avdd.n439 avdd.n112 16.3134
R7290 avdd.n81 avdd.n79 15.7779
R7291 avdd.n19 avdd.n18 15.5799
R7292 avdd.n18 avdd.n0 15.5799
R7293 avdd.n31 avdd.n30 15.5799
R7294 avdd.n187 avdd.n185 15.4172
R7295 avdd.n193 avdd.n185 15.4172
R7296 avdd.n183 avdd.n176 15.4172
R7297 avdd.n184 avdd.n183 15.4172
R7298 avdd.n179 avdd.n177 15.4172
R7299 avdd.n190 avdd.n186 15.4172
R7300 avdd.n386 avdd.t98 13.848
R7301 avdd.n386 avdd.t85 13.848
R7302 avdd.n388 avdd.t5 13.848
R7303 avdd.n388 avdd.t101 13.848
R7304 avdd.n390 avdd.t83 13.848
R7305 avdd.n390 avdd.t87 13.848
R7306 avdd.n531 avdd.n530 13.5116
R7307 avdd.n79 avdd.n78 13.3823
R7308 avdd.n506 avdd.n474 13.2339
R7309 avdd.n501 avdd.n500 13.2148
R7310 avdd.n501 avdd.t20 13.2148
R7311 avdd.n519 avdd.n518 13.2148
R7312 avdd.n519 avdd.t20 13.2148
R7313 avdd.n468 avdd.n461 13.2148
R7314 avdd.n511 avdd.n477 13.2148
R7315 avdd.n477 avdd.t20 13.2148
R7316 avdd.n466 avdd.n460 13.2148
R7317 avdd.t116 avdd.n466 13.2148
R7318 avdd.n490 avdd.n489 13.2148
R7319 avdd.t118 avdd.n490 13.2148
R7320 avdd.n495 avdd.n467 13.2148
R7321 avdd.t116 avdd.n467 13.2148
R7322 avdd.n484 avdd.n478 13.2148
R7323 avdd.n107 avdd.n106 13.0717
R7324 avdd.n531 avdd.n462 12.9974
R7325 avdd.n79 avdd.n53 12.4253
R7326 avdd.n46 avdd.n35 12.3338
R7327 avdd.n46 avdd.n40 12.3338
R7328 avdd.n105 avdd.n104 12.3338
R7329 avdd.n104 avdd.n103 12.3338
R7330 avdd.n100 avdd.n97 12.3338
R7331 avdd.n85 avdd.n44 12.3338
R7332 avdd.n45 avdd.n44 12.3338
R7333 avdd.n430 avdd.t113 12.1529
R7334 avdd.n93 avdd.n92 11.2161
R7335 avdd.n94 avdd.n36 11.2161
R7336 avdd.n32 avdd.n31 10.8988
R7337 avdd.n81 avdd.n80 10.809
R7338 avdd.n465 avdd.n462 9.99435
R7339 avdd.n442 avdd.n438 9.70387
R7340 avdd.n443 avdd.n113 9.61683
R7341 avdd.n125 avdd.t89 9.5505
R7342 avdd.n125 avdd.t91 9.5505
R7343 avdd.n126 avdd.t1 9.5505
R7344 avdd.n126 avdd.t3 9.5505
R7345 avdd.n127 avdd.t81 9.5505
R7346 avdd.n127 avdd.t22 9.5505
R7347 avdd.n92 avdd.n43 9.55042
R7348 avdd.n279 avdd.n278 9.3395
R7349 avdd.n280 avdd.n279 9.3005
R7350 avdd.n282 avdd.n280 9.3005
R7351 avdd.n282 avdd.n281 9.3005
R7352 avdd.n281 avdd.n279 9.3005
R7353 avdd.n296 avdd.n294 9.3005
R7354 avdd.n313 avdd.n263 9.3005
R7355 avdd.n265 avdd.n263 9.3005
R7356 avdd.n311 avdd.n263 9.3005
R7357 avdd.n317 avdd.n256 9.3005
R7358 avdd.n321 avdd.n317 9.3005
R7359 avdd.n317 avdd.n315 9.3005
R7360 avdd.n335 avdd.n244 9.3005
R7361 avdd.n244 avdd.n242 9.3005
R7362 avdd.n333 avdd.n244 9.3005
R7363 avdd.n252 avdd.n246 9.3005
R7364 avdd.n373 avdd.n223 9.3005
R7365 avdd.n375 avdd.n223 9.3005
R7366 avdd.n223 avdd.n221 9.3005
R7367 avdd.n366 avdd.n231 9.3005
R7368 avdd.n368 avdd.n231 9.3005
R7369 avdd.n231 avdd.n226 9.3005
R7370 avdd.n360 avdd.n358 9.3005
R7371 avdd.n358 avdd.n357 9.3005
R7372 avdd.n298 avdd.n297 9.3005
R7373 avdd.n297 avdd.n296 9.3005
R7374 avdd.n297 avdd.n274 9.3005
R7375 avdd.n313 avdd.n312 9.3005
R7376 avdd.n312 avdd.n311 9.3005
R7377 avdd.n312 avdd.n265 9.3005
R7378 avdd.n320 avdd.n256 9.3005
R7379 avdd.n320 avdd.n315 9.3005
R7380 avdd.n321 avdd.n320 9.3005
R7381 avdd.n335 avdd.n334 9.3005
R7382 avdd.n334 avdd.n333 9.3005
R7383 avdd.n334 avdd.n242 9.3005
R7384 avdd.n251 avdd.n214 9.3005
R7385 avdd.n252 avdd.n251 9.3005
R7386 avdd.n251 avdd.n250 9.3005
R7387 avdd.n374 avdd.n373 9.3005
R7388 avdd.n374 avdd.n221 9.3005
R7389 avdd.n375 avdd.n374 9.3005
R7390 avdd.n367 avdd.n366 9.3005
R7391 avdd.n367 avdd.n226 9.3005
R7392 avdd.n368 avdd.n367 9.3005
R7393 avdd.n359 avdd.n357 9.3005
R7394 avdd.n360 avdd.n359 9.3005
R7395 avdd.n284 avdd.n283 9.3005
R7396 avdd.n276 avdd.n275 9.3005
R7397 avdd.n292 avdd.n291 9.3005
R7398 avdd.n295 avdd.n271 9.3005
R7399 avdd.n300 avdd.n299 9.3005
R7400 avdd.n267 avdd.n266 9.3005
R7401 avdd.n310 avdd.n309 9.3005
R7402 avdd.n308 avdd.n261 9.3005
R7403 avdd.n314 avdd.n260 9.3005
R7404 avdd.n323 avdd.n322 9.3005
R7405 avdd.n318 avdd.n257 9.3005
R7406 avdd.n331 avdd.n330 9.3005
R7407 avdd.n332 avdd.n240 9.3005
R7408 avdd.n337 avdd.n336 9.3005
R7409 avdd.n254 avdd.n241 9.3005
R7410 avdd.n253 avdd.n238 9.3005
R7411 avdd.n247 avdd.n216 9.3005
R7412 avdd.n380 avdd.n379 9.3005
R7413 avdd.n378 avdd.n215 9.3005
R7414 avdd.n377 avdd.n376 9.3005
R7415 avdd.n224 avdd.n220 9.3005
R7416 avdd.n372 avdd.n371 9.3005
R7417 avdd.n370 avdd.n369 9.3005
R7418 avdd.n232 avdd.n229 9.3005
R7419 avdd.n365 avdd.n364 9.3005
R7420 avdd.n363 avdd.n234 9.3005
R7421 avdd.n362 avdd.n361 9.3005
R7422 avdd.n472 avdd.n468 9.21551
R7423 avdd.n485 avdd.n484 9.21551
R7424 avdd.n327 avdd.t66 8.69615
R7425 avdd.t48 avdd.n355 8.69615
R7426 avdd.t13 avdd.n28 7.23338
R7427 avdd.t14 avdd.n12 7.23338
R7428 avdd.n408 avdd.n398 6.85235
R7429 avdd.n430 avdd.n398 6.85235
R7430 avdd.n432 avdd.n431 6.85235
R7431 avdd.n431 avdd.n430 6.85235
R7432 avdd.n526 avdd.n525 6.79556
R7433 avdd.n437 avdd 6.67576
R7434 avdd.n530 avdd.n463 6.63754
R7435 avdd.n124 avdd.n123 6.60764
R7436 avdd.n123 avdd.n122 6.60764
R7437 avdd.n440 avdd.n115 6.56673
R7438 avdd.n441 avdd.n124 6.56673
R7439 avdd.n94 avdd.n93 6.54643
R7440 avdd.n101 avdd.n36 6.54643
R7441 avdd.n65 avdd.n64 5.85127
R7442 avdd.n413 avdd.t6 5.81251
R7443 avdd.n443 avdd.n442 5.42014
R7444 avdd.n433 avdd.n432 5.33383
R7445 avdd.n532 avdd.n460 5.19808
R7446 avdd.n69 avdd.n68 4.97214
R7447 avdd.n67 avdd.n54 4.88297
R7448 avdd.n471 avdd.n465 4.87435
R7449 avdd.n508 avdd.n474 4.76501
R7450 avdd.n32 avdd.n0 4.68164
R7451 avdd.n72 avdd.n71 4.67841
R7452 avdd.n528 avdd.n527 4.67518
R7453 avdd.n294 avdd.n272 4.64202
R7454 avdd.n249 avdd.n246 4.64202
R7455 avdd.n527 avdd.n463 4.43127
R7456 avdd.n77 avdd.n56 4.41262
R7457 avdd.n455 avdd.n114 4.36414
R7458 avdd.t55 avdd.n269 4.34833
R7459 avdd.n345 avdd.t64 4.34833
R7460 avdd.n85 avdd.n34 4.20442
R7461 avdd.t111 avdd.n96 4.16651
R7462 avdd.n212 avdd.t120 4.16123
R7463 avdd.t118 avdd.n485 3.92667
R7464 avdd.n472 avdd.t20 3.92667
R7465 avdd.n439 avdd.n438 3.83483
R7466 avdd.n445 avdd.n444 3.15894
R7467 avdd.n509 avdd.n508 3.12119
R7468 avdd.n78 avdd.n54 3.0725
R7469 avdd.n64 avdd.n43 3.01226
R7470 avdd.n528 avdd.n464 2.85313
R7471 avdd.n382 avdd.n381 2.64322
R7472 avdd.n436 avdd.n384 2.63743
R7473 avdd.n435 avdd.n434 2.59863
R7474 avdd.n479 avdd 2.5005
R7475 avdd.n69 avdd.n59 2.47792
R7476 avdd.n170 avdd.n169 2.41559
R7477 avdd.n493 avdd.n481 2.36947
R7478 avdd.n530 avdd.n529 2.3255
R7479 avdd.n145 avdd.n133 2.17789
R7480 avdd.n66 avdd.n65 2.10699
R7481 avdd.n86 avdd.n43 2.07109
R7482 avdd.n536 avdd.n111 1.86784
R7483 avdd.n453 avdd.n452 1.72947
R7484 avdd.n452 avdd.n451 1.72947
R7485 avdd.n509 avdd.n464 1.66013
R7486 avdd.n213 avdd.n212 1.46404
R7487 avdd.n148 avdd.n145 1.44956
R7488 avdd.n536 avdd.n535 1.43719
R7489 avdd.n445 avdd.n120 1.3811
R7490 avdd.n121 avdd.n120 1.3811
R7491 avdd.n437 avdd.n436 1.37352
R7492 avdd.n448 avdd.n447 1.36079
R7493 avdd.n449 avdd.n448 1.36079
R7494 avdd.n107 avdd.n105 1.30227
R7495 avdd.n109 avdd.n34 1.30044
R7496 avdd.n108 avdd.n35 1.30044
R7497 avdd.n507 avdd.n506 1.21911
R7498 avdd.n171 avdd.n133 1.19205
R7499 avdd.n172 avdd.n171 1.1255
R7500 avdd.n458 avdd.n457 1.1255
R7501 avdd.n535 avdd.n458 0.998081
R7502 avdd.n497 avdd.n471 0.985115
R7503 avdd.n481 avdd.n480 0.974799
R7504 avdd.n171 avdd.n170 0.97298
R7505 avdd.n384 avdd.n382 0.959959
R7506 avdd.n80 avdd.n43 0.951668
R7507 avdd.n86 avdd.n85 0.847559
R7508 avdd.n384 avdd.n383 0.844173
R7509 avdd.n158 avdd.n157 0.839844
R7510 avdd.n208 avdd.n175 0.780195
R7511 avdd.n435 avdd.n385 0.742984
R7512 avdd.n525 avdd.n463 0.711611
R7513 avdd.n68 avdd.n63 0.657216
R7514 avdd.n510 avdd.n509 0.6205
R7515 avdd.n537 avdd.n32 0.610562
R7516 avdd.n447 avdd.n446 0.565206
R7517 avdd.n209 avdd.n208 0.554667
R7518 avdd.n385 avdd.t122 0.545513
R7519 avdd.n537 avdd.n536 0.532487
R7520 avdd.n434 avdd.n393 0.525114
R7521 avdd.n116 avdd.n115 0.496479
R7522 avdd.n118 avdd.n116 0.496479
R7523 avdd.n434 avdd.n433 0.464249
R7524 avdd.n157 avdd.n133 0.404848
R7525 avdd.n117 avdd.n114 0.363958
R7526 avdd.n450 avdd.n117 0.363958
R7527 avdd.n382 avdd.n213 0.35824
R7528 avdd.n507 avdd.n459 0.354021
R7529 avdd.n498 avdd.n464 0.344944
R7530 avdd.n442 avdd.n441 0.344944
R7531 avdd.n62 avdd.n61 0.319135
R7532 avdd.n389 avdd.n387 0.316214
R7533 avdd.n392 avdd.n391 0.312643
R7534 avdd.n391 avdd.n389 0.312643
R7535 avdd.n72 avdd.n59 0.308934
R7536 avdd.n78 avdd.n77 0.291409
R7537 avdd.n67 avdd.n66 0.271595
R7538 avdd.n173 avdd.n172 0.266737
R7539 avdd.n56 avdd.n55 0.248242
R7540 avdd.n80 avdd.n33 0.238962
R7541 avdd.n62 avdd.n60 0.237956
R7542 avdd avdd.n537 0.236316
R7543 avdd.n383 avdd.t25 0.232449
R7544 avdd.n383 avdd.t121 0.231345
R7545 avdd.n480 avdd 0.22534
R7546 avdd.n436 avdd.n435 0.209118
R7547 avdd.n63 avdd.n60 0.202509
R7548 avdd.n457 avdd.n112 0.200606
R7549 avdd avdd.n392 0.199071
R7550 avdd.n533 avdd.n532 0.190296
R7551 avdd.n174 avdd.n173 0.182805
R7552 avdd.n210 avdd.n209 0.180916
R7553 avdd.n212 avdd.n211 0.174607
R7554 avdd.n108 avdd.n107 0.17436
R7555 avdd.n109 avdd.n108 0.173953
R7556 avdd.n454 avdd.n453 0.159506
R7557 avdd.n458 avdd 0.133565
R7558 avdd.n534 avdd 0.123304
R7559 avdd.n446 avdd.n113 0.115323
R7560 avdd.n533 avdd.n459 0.102337
R7561 avdd.n211 avdd.n210 0.100311
R7562 avdd.n511 avdd.n510 0.0989615
R7563 avdd.n454 avdd.n112 0.0969049
R7564 avdd.n130 avdd.n129 0.0771667
R7565 avdd.n479 avdd 0.0758012
R7566 avdd.n132 avdd.n131 0.0757381
R7567 avdd.n444 avdd.n443 0.0743095
R7568 avdd.n385 avdd.t99 0.0677395
R7569 avdd.n129 avdd.n128 0.0650238
R7570 avdd.n131 avdd.n130 0.0633571
R7571 avdd.n529 avdd.n459 0.060719
R7572 avdd.n508 avdd.n507 0.0567495
R7573 avdd.n68 avdd.n67 0.0485456
R7574 avdd.n292 avdd.n275 0.0485
R7575 avdd.n299 avdd.n266 0.0485
R7576 avdd.n332 avdd.n331 0.0485
R7577 avdd.n254 avdd.n253 0.0485
R7578 avdd.n380 avdd.n215 0.0485
R7579 avdd.n365 avdd.n234 0.0485
R7580 avdd.n110 avdd.n109 0.0448811
R7581 avdd.n315 avdd.n314 0.044
R7582 avdd.n372 avdd.n226 0.044
R7583 avdd.n314 avdd.n313 0.041
R7584 avdd.n373 avdd.n372 0.041
R7585 avdd.n66 avdd.n33 0.0404023
R7586 avdd.n438 avdd.n437 0.0362143
R7587 avdd.n393 avdd 0.0355
R7588 avdd.n111 avdd.n110 0.0345909
R7589 avdd avdd.n111 0.0339677
R7590 avdd.n361 avdd.n357 0.0335
R7591 avdd.n110 avdd.n33 0.0326661
R7592 avdd.n172 avdd.n132 0.0324048
R7593 avdd.n311 avdd.n266 0.032
R7594 avdd.n322 avdd.n321 0.032
R7595 avdd.n336 avdd.n335 0.032
R7596 avdd.n221 avdd.n215 0.032
R7597 avdd.n369 avdd.n368 0.032
R7598 avdd.n296 avdd.n295 0.029
R7599 avdd.n265 avdd.n261 0.029
R7600 avdd.n331 avdd.n256 0.029
R7601 avdd.n252 avdd.n247 0.029
R7602 avdd.n375 avdd.n224 0.029
R7603 avdd.n366 avdd.n365 0.029
R7604 avdd.n529 avdd.n528 0.0287623
R7605 avdd.n283 avdd.n282 0.0275
R7606 avdd.n535 avdd.n534 0.0272857
R7607 avdd.n440 avdd.n439 0.0267712
R7608 avdd.n282 avdd.n275 0.0215
R7609 avdd.n360 avdd 0.0215
R7610 avdd.n296 avdd.n292 0.02
R7611 avdd.n310 avdd.n265 0.02
R7612 avdd.n318 avdd.n256 0.02
R7613 avdd avdd.n242 0.02
R7614 avdd.n253 avdd.n252 0.02
R7615 avdd.n376 avdd.n375 0.02
R7616 avdd.n366 avdd.n232 0.02
R7617 avdd.n456 avdd.n455 0.0199154
R7618 avdd.n274 avdd.n272 0.0189652
R7619 avdd.n250 avdd.n249 0.0189652
R7620 avdd.n298 avdd.n272 0.0189652
R7621 avdd.n249 avdd.n214 0.0189652
R7622 avdd.n480 avdd 0.0182716
R7623 avdd.n311 avdd.n310 0.017
R7624 avdd.n321 avdd.n318 0.017
R7625 avdd.n333 avdd 0.017
R7626 avdd.n335 avdd.n254 0.017
R7627 avdd.n376 avdd.n221 0.017
R7628 avdd.n368 avdd.n232 0.017
R7629 avdd.n357 avdd.n234 0.0155
R7630 avdd.n534 avdd.n533 0.0118818
R7631 avdd.n211 avdd 0.0105756
R7632 avdd.n283 avdd.n279 0.0095
R7633 avdd.n209 avdd.n174 0.00805668
R7634 avdd.n295 avdd.n274 0.008
R7635 avdd.n313 avdd.n261 0.008
R7636 avdd.n333 avdd.n332 0.008
R7637 avdd.n250 avdd.n247 0.008
R7638 avdd.n373 avdd.n224 0.008
R7639 avdd avdd.n479 0.00629073
R7640 avdd.n299 avdd.n298 0.005
R7641 avdd.n322 avdd.n315 0.005
R7642 avdd.n336 avdd.n242 0.005
R7643 avdd.n369 avdd.n226 0.005
R7644 avdd.n213 avdd 0.00364861
R7645 avdd.n381 avdd.n380 0.0035
R7646 avdd.n361 avdd.n360 0.0035
R7647 avdd.n381 avdd.n214 0.002
R7648 a_25251_n288267.n2 a_25251_n288267.t3 341.087
R7649 a_25251_n288267.t1 a_25251_n288267.n2 340.214
R7650 a_25251_n288267.n2 a_25251_n288267.t2 232.124
R7651 a_25251_n288267.n1 a_25251_n288267.t5 173.871
R7652 a_25251_n288267.n0 a_25251_n288267.t4 173.868
R7653 a_25251_n288267.n1 a_25251_n288267.t6 164.47
R7654 a_25251_n288267.n0 a_25251_n288267.t0 4.32892
R7655 a_25251_n288267.n2 a_25251_n288267.n1 3.0715
R7656 a_25251_n288267.n1 a_25251_n288267.n0 2.23288
R7657 a_25567_n288267.t3 a_25567_n288267.n1 341.103
R7658 a_25567_n288267.n1 a_25567_n288267.t2 340.214
R7659 a_25567_n288267.n1 a_25567_n288267.t1 232.145
R7660 a_25567_n288267.n0 a_25567_n288267.t6 175.047
R7661 a_25567_n288267.n0 a_25567_n288267.t4 173.871
R7662 a_25567_n288267.n0 a_25567_n288267.t5 164.475
R7663 a_25567_n288267.n1 a_25567_n288267.t0 6.76699
R7664 a_25567_n288267.n1 a_25567_n288267.n0 3.77356
R7665 porb_h[1].n2 porb_h[1].n1 157.593
R7666 porb_h[1].n8 porb_h[1].n7 157.591
R7667 porb_h[1].n12 porb_h[1].n11 157.591
R7668 porb_h[1].n16 porb_h[1].n15 157.591
R7669 porb_h[1].n20 porb_h[1].n19 157.591
R7670 porb_h[1].n24 porb_h[1].n23 157.591
R7671 porb_h[1].n28 porb_h[1].n27 157.591
R7672 porb_h[1].n32 porb_h[1].n31 157.591
R7673 porb_h[1].n8 porb_h[1].n6 136.965
R7674 porb_h[1].n12 porb_h[1].n10 136.965
R7675 porb_h[1].n16 porb_h[1].n14 136.965
R7676 porb_h[1].n20 porb_h[1].n18 136.965
R7677 porb_h[1].n24 porb_h[1].n22 136.965
R7678 porb_h[1].n28 porb_h[1].n26 136.965
R7679 porb_h[1].n32 porb_h[1].n30 136.965
R7680 porb_h[1].n2 porb_h[1].n0 136.965
R7681 porb_h[1].n6 porb_h[1].t0 21.2805
R7682 porb_h[1].n6 porb_h[1].t15 21.2805
R7683 porb_h[1].n10 porb_h[1].t11 21.2805
R7684 porb_h[1].n10 porb_h[1].t5 21.2805
R7685 porb_h[1].n14 porb_h[1].t12 21.2805
R7686 porb_h[1].n14 porb_h[1].t4 21.2805
R7687 porb_h[1].n18 porb_h[1].t7 21.2805
R7688 porb_h[1].n18 porb_h[1].t13 21.2805
R7689 porb_h[1].n22 porb_h[1].t14 21.2805
R7690 porb_h[1].n22 porb_h[1].t8 21.2805
R7691 porb_h[1].n26 porb_h[1].t10 21.2805
R7692 porb_h[1].n26 porb_h[1].t2 21.2805
R7693 porb_h[1].n30 porb_h[1].t3 21.2805
R7694 porb_h[1].n30 porb_h[1].t1 21.2805
R7695 porb_h[1].n0 porb_h[1].t9 21.2805
R7696 porb_h[1].n0 porb_h[1].t6 21.2805
R7697 porb_h[1].n7 porb_h[1].t29 17.8272
R7698 porb_h[1].n7 porb_h[1].t28 17.8272
R7699 porb_h[1].n11 porb_h[1].t25 17.8272
R7700 porb_h[1].n11 porb_h[1].t17 17.8272
R7701 porb_h[1].n15 porb_h[1].t24 17.8272
R7702 porb_h[1].n15 porb_h[1].t16 17.8272
R7703 porb_h[1].n19 porb_h[1].t19 17.8272
R7704 porb_h[1].n19 porb_h[1].t26 17.8272
R7705 porb_h[1].n23 porb_h[1].t27 17.8272
R7706 porb_h[1].n23 porb_h[1].t22 17.8272
R7707 porb_h[1].n27 porb_h[1].t23 17.8272
R7708 porb_h[1].n27 porb_h[1].t31 17.8272
R7709 porb_h[1].n31 porb_h[1].t18 17.8272
R7710 porb_h[1].n31 porb_h[1].t30 17.8272
R7711 porb_h[1].n1 porb_h[1].t21 17.8272
R7712 porb_h[1].n1 porb_h[1].t20 17.8272
R7713 porb_h[1].n3 porb_h[1].n2 9.98018
R7714 porb_h[1].n9 porb_h[1].n8 9.98018
R7715 porb_h[1].n13 porb_h[1].n12 9.98018
R7716 porb_h[1].n17 porb_h[1].n16 9.98018
R7717 porb_h[1].n21 porb_h[1].n20 9.98018
R7718 porb_h[1].n25 porb_h[1].n24 9.98018
R7719 porb_h[1].n29 porb_h[1].n28 9.98018
R7720 porb_h[1].n33 porb_h[1].n32 9.98018
R7721 porb_h[1].n34 porb_h[1].n33 2.13429
R7722 porb_h[1].n35 porb_h[1] 1.4032
R7723 porb_h[1].n33 porb_h[1].n29 0.379141
R7724 porb_h[1].n29 porb_h[1].n25 0.379141
R7725 porb_h[1].n25 porb_h[1].n21 0.379141
R7726 porb_h[1].n21 porb_h[1].n17 0.379141
R7727 porb_h[1].n17 porb_h[1].n13 0.379141
R7728 porb_h[1].n13 porb_h[1].n9 0.379141
R7729 porb_h[1].n9 porb_h[1].n5 0.28084
R7730 porb_h[1].n4 porb_h[1] 0.213735
R7731 porb_h[1].n5 porb_h[1].n4 0.191676
R7732 porb_h[1].n34 porb_h[1] 0.186724
R7733 porb_h[1].n5 porb_h[1] 0.133995
R7734 porb_h[1].n4 porb_h[1].n3 0.0793043
R7735 porb_h[1].n3 porb_h[1] 0.0793043
R7736 porb_h[1].n35 porb_h[1].n34 0.0693775
R7737 porb_h[1] porb_h[1].n35 0.0305245
R7738 a_34073_n287091.t5 a_34073_n287091.n0 166.194
R7739 a_34073_n287091.n4 a_34073_n287091.n0 1.67896
R7740 a_34073_n287091.t6 a_34073_n287091.n6 332.308
R7741 a_34073_n287091.t9 a_34073_n287091.n0 165.965
R7742 a_34073_n287091.t7 a_34073_n287091.n3 331.928
R7743 a_34073_n287091.n6 a_34073_n287091.t7 331.928
R7744 a_34073_n287091.n3 a_34073_n287091.t6 331.928
R7745 a_34073_n287091.n4 a_34073_n287091.t8 138.482
R7746 a_34073_n287091.n1 a_34073_n287091.t1 86.002
R7747 a_34073_n287091.n1 a_34073_n287091.t0 85.9222
R7748 a_34073_n287091.n1 a_34073_n287091.t2 49.8929
R7749 a_34073_n287091.t3 a_34073_n287091.n1 49.8725
R7750 a_34073_n287091.n5 a_34073_n287091.t4 4.72862
R7751 a_34073_n287091.n2 a_34073_n287091.n4 0.323471
R7752 a_34073_n287091.n2 a_34073_n287091.n1 1.06604
R7753 a_34073_n287091.n6 a_34073_n287091.n5 1.84029
R7754 a_34073_n287091.n5 a_34073_n287091.n3 1.06414
R7755 a_34073_n287091.n2 a_34073_n287091.n3 1.63985
R7756 a_35454_n291454.t28 a_35454_n291454.t39 353.467
R7757 a_35454_n291454.t49 a_35454_n291454.t59 353.467
R7758 a_35454_n291454.t63 a_35454_n291454.t27 353.467
R7759 a_35454_n291454.t37 a_35454_n291454.t48 353.467
R7760 a_35454_n291454.t53 a_35454_n291454.t62 353.467
R7761 a_35454_n291454.t24 a_35454_n291454.t36 353.467
R7762 a_35454_n291454.t46 a_35454_n291454.t57 353.467
R7763 a_35454_n291454.t34 a_35454_n291454.t44 353.467
R7764 a_35454_n291454.t55 a_35454_n291454.t64 353.467
R7765 a_35454_n291454.t69 a_35454_n291454.t32 353.467
R7766 a_35454_n291454.t42 a_35454_n291454.t54 353.467
R7767 a_35454_n291454.t61 a_35454_n291454.t25 353.467
R7768 a_35454_n291454.t30 a_35454_n291454.t41 353.467
R7769 a_35454_n291454.t51 a_35454_n291454.t60 353.467
R7770 a_35454_n291454.t66 a_35454_n291454.t29 353.467
R7771 a_35454_n291454.t38 a_35454_n291454.t50 353.467
R7772 a_35454_n291454.n12 a_35454_n291454.n10 299.851
R7773 a_35454_n291454.n8 a_35454_n291454.n6 299.851
R7774 a_35454_n291454.n4 a_35454_n291454.n2 299.851
R7775 a_35454_n291454.n50 a_35454_n291454.n49 299.851
R7776 a_35454_n291454.n49 a_35454_n291454.n48 299.414
R7777 a_35454_n291454.n12 a_35454_n291454.n11 299.414
R7778 a_35454_n291454.n8 a_35454_n291454.n7 299.414
R7779 a_35454_n291454.n4 a_35454_n291454.n3 299.414
R7780 a_35454_n291454.n14 a_35454_n291454.t28 232.382
R7781 a_35454_n291454.n21 a_35454_n291454.t38 232.382
R7782 a_35454_n291454.n47 a_35454_n291454.n1 197.123
R7783 a_35454_n291454.n0 a_35454_n291454.n13 197.123
R7784 a_35454_n291454.n45 a_35454_n291454.n9 197.123
R7785 a_35454_n291454.n46 a_35454_n291454.n5 197.123
R7786 a_35454_n291454.n36 a_35454_n291454.t33 185.79
R7787 a_35454_n291454.n29 a_35454_n291454.t70 185.79
R7788 a_35454_n291454.n14 a_35454_n291454.t49 162.274
R7789 a_35454_n291454.n15 a_35454_n291454.t63 162.274
R7790 a_35454_n291454.n16 a_35454_n291454.t37 162.274
R7791 a_35454_n291454.n17 a_35454_n291454.t53 162.274
R7792 a_35454_n291454.n18 a_35454_n291454.t24 162.274
R7793 a_35454_n291454.n19 a_35454_n291454.t46 162.274
R7794 a_35454_n291454.n20 a_35454_n291454.t34 162.274
R7795 a_35454_n291454.n27 a_35454_n291454.t55 162.274
R7796 a_35454_n291454.n26 a_35454_n291454.t69 162.274
R7797 a_35454_n291454.n25 a_35454_n291454.t42 162.274
R7798 a_35454_n291454.n24 a_35454_n291454.t61 162.274
R7799 a_35454_n291454.n23 a_35454_n291454.t30 162.274
R7800 a_35454_n291454.n22 a_35454_n291454.t51 162.274
R7801 a_35454_n291454.n21 a_35454_n291454.t66 162.274
R7802 a_35454_n291454.n36 a_35454_n291454.t65 115.68
R7803 a_35454_n291454.n37 a_35454_n291454.t45 115.68
R7804 a_35454_n291454.n38 a_35454_n291454.t71 115.68
R7805 a_35454_n291454.n39 a_35454_n291454.t56 115.68
R7806 a_35454_n291454.n40 a_35454_n291454.t35 115.68
R7807 a_35454_n291454.n41 a_35454_n291454.t68 115.68
R7808 a_35454_n291454.n42 a_35454_n291454.t47 115.68
R7809 a_35454_n291454.n35 a_35454_n291454.t26 115.68
R7810 a_35454_n291454.n34 a_35454_n291454.t40 115.68
R7811 a_35454_n291454.n33 a_35454_n291454.t67 115.68
R7812 a_35454_n291454.n32 a_35454_n291454.t52 115.68
R7813 a_35454_n291454.n31 a_35454_n291454.t31 115.68
R7814 a_35454_n291454.n30 a_35454_n291454.t58 115.68
R7815 a_35454_n291454.n29 a_35454_n291454.t43 115.68
R7816 a_35454_n291454.n30 a_35454_n291454.n29 70.1096
R7817 a_35454_n291454.n31 a_35454_n291454.n30 70.1096
R7818 a_35454_n291454.n32 a_35454_n291454.n31 70.1096
R7819 a_35454_n291454.n33 a_35454_n291454.n32 70.1096
R7820 a_35454_n291454.n34 a_35454_n291454.n33 70.1096
R7821 a_35454_n291454.n35 a_35454_n291454.n34 70.1096
R7822 a_35454_n291454.n42 a_35454_n291454.n41 70.1096
R7823 a_35454_n291454.n41 a_35454_n291454.n40 70.1096
R7824 a_35454_n291454.n40 a_35454_n291454.n39 70.1096
R7825 a_35454_n291454.n39 a_35454_n291454.n38 70.1096
R7826 a_35454_n291454.n38 a_35454_n291454.n37 70.1096
R7827 a_35454_n291454.n37 a_35454_n291454.n36 70.1096
R7828 a_35454_n291454.n15 a_35454_n291454.n14 70.1096
R7829 a_35454_n291454.n16 a_35454_n291454.n15 70.1096
R7830 a_35454_n291454.n17 a_35454_n291454.n16 70.1096
R7831 a_35454_n291454.n18 a_35454_n291454.n17 70.1096
R7832 a_35454_n291454.n19 a_35454_n291454.n18 70.1096
R7833 a_35454_n291454.n20 a_35454_n291454.n19 70.1096
R7834 a_35454_n291454.n27 a_35454_n291454.n26 70.1096
R7835 a_35454_n291454.n26 a_35454_n291454.n25 70.1096
R7836 a_35454_n291454.n25 a_35454_n291454.n24 70.1096
R7837 a_35454_n291454.n24 a_35454_n291454.n23 70.1096
R7838 a_35454_n291454.n23 a_35454_n291454.n22 70.1096
R7839 a_35454_n291454.n22 a_35454_n291454.n21 70.1096
R7840 a_35454_n291454.n48 a_35454_n291454.t10 46.4362
R7841 a_35454_n291454.n48 a_35454_n291454.t21 46.4362
R7842 a_35454_n291454.n10 a_35454_n291454.t8 46.4362
R7843 a_35454_n291454.n10 a_35454_n291454.t13 46.4362
R7844 a_35454_n291454.n11 a_35454_n291454.t12 46.4362
R7845 a_35454_n291454.n11 a_35454_n291454.t18 46.4362
R7846 a_35454_n291454.n6 a_35454_n291454.t15 46.4362
R7847 a_35454_n291454.n6 a_35454_n291454.t9 46.4362
R7848 a_35454_n291454.n7 a_35454_n291454.t19 46.4362
R7849 a_35454_n291454.n7 a_35454_n291454.t14 46.4362
R7850 a_35454_n291454.n2 a_35454_n291454.t20 46.4362
R7851 a_35454_n291454.n2 a_35454_n291454.t11 46.4362
R7852 a_35454_n291454.n3 a_35454_n291454.t22 46.4362
R7853 a_35454_n291454.n3 a_35454_n291454.t16 46.4362
R7854 a_35454_n291454.t23 a_35454_n291454.n50 46.4362
R7855 a_35454_n291454.n50 a_35454_n291454.t17 46.4362
R7856 a_35454_n291454.n1 a_35454_n291454.t1 39.6005
R7857 a_35454_n291454.n1 a_35454_n291454.t7 39.6005
R7858 a_35454_n291454.n13 a_35454_n291454.t3 39.6005
R7859 a_35454_n291454.n13 a_35454_n291454.t5 39.6005
R7860 a_35454_n291454.n9 a_35454_n291454.t6 39.6005
R7861 a_35454_n291454.n9 a_35454_n291454.t2 39.6005
R7862 a_35454_n291454.n5 a_35454_n291454.t0 39.6005
R7863 a_35454_n291454.n5 a_35454_n291454.t4 39.6005
R7864 a_35454_n291454.n43 a_35454_n291454.n35 35.055
R7865 a_35454_n291454.n43 a_35454_n291454.n42 35.055
R7866 a_35454_n291454.n28 a_35454_n291454.n20 35.055
R7867 a_35454_n291454.n28 a_35454_n291454.n27 35.055
R7868 a_35454_n291454.n44 a_35454_n291454.n43 10.2069
R7869 a_35454_n291454.n44 a_35454_n291454.n28 10.156
R7870 a_35454_n291454.n0 a_35454_n291454.n44 2.6231
R7871 a_35454_n291454.n0 a_35454_n291454.n12 0.504406
R7872 a_35454_n291454.n45 a_35454_n291454.n8 0.504406
R7873 a_35454_n291454.n46 a_35454_n291454.n4 0.504406
R7874 a_35454_n291454.n49 a_35454_n291454.n47 0.504406
R7875 a_35454_n291454.n46 a_35454_n291454.n45 0.276362
R7876 a_35454_n291454.n47 a_35454_n291454.n46 0.276362
R7877 a_35454_n291454.n45 a_35454_n291454.n0 0.276362
R7878 por.n6 por.n4 299.851
R7879 por.n10 por.n8 299.851
R7880 por.n14 por.n12 299.851
R7881 por.n18 por.n16 299.851
R7882 por.n22 por.n20 299.851
R7883 por.n26 por.n24 299.851
R7884 por.n30 por.n28 299.851
R7885 por.n2 por.n0 299.851
R7886 por.n6 por.n5 299.414
R7887 por.n10 por.n9 299.414
R7888 por.n14 por.n13 299.414
R7889 por.n18 por.n17 299.414
R7890 por.n22 por.n21 299.414
R7891 por.n26 por.n25 299.414
R7892 por.n30 por.n29 299.414
R7893 por.n2 por.n1 299.414
R7894 por.n38 por.n7 197.123
R7895 por.n37 por.n11 197.123
R7896 por.n36 por.n15 197.123
R7897 por.n35 por.n19 197.123
R7898 por.n34 por.n23 197.123
R7899 por.n33 por.n27 197.123
R7900 por.n32 por.n31 197.123
R7901 por.n39 por.n3 197.094
R7902 por.n4 por.t45 46.4362
R7903 por.n4 por.t31 46.4362
R7904 por.n5 por.t19 46.4362
R7905 por.n5 por.t38 46.4362
R7906 por.n8 por.t20 46.4362
R7907 por.n8 por.t39 46.4362
R7908 por.n9 por.t27 46.4362
R7909 por.n9 por.t47 46.4362
R7910 por.n12 por.t24 46.4362
R7911 por.n12 por.t33 46.4362
R7912 por.n13 por.t32 46.4362
R7913 por.n13 por.t40 46.4362
R7914 por.n16 por.t18 46.4362
R7915 por.n16 por.t41 46.4362
R7916 por.n17 por.t25 46.4362
R7917 por.n17 por.t16 46.4362
R7918 por.n20 por.t26 46.4362
R7919 por.n20 por.t46 46.4362
R7920 por.n21 por.t34 46.4362
R7921 por.n21 por.t21 46.4362
R7922 por.n24 por.t35 46.4362
R7923 por.n24 por.t22 46.4362
R7924 por.n25 por.t42 46.4362
R7925 por.n25 por.t28 46.4362
R7926 por.n28 por.t43 46.4362
R7927 por.n28 por.t29 46.4362
R7928 por.n29 por.t17 46.4362
R7929 por.n29 por.t37 46.4362
R7930 por.n0 por.t36 46.4362
R7931 por.n0 por.t23 46.4362
R7932 por.n1 por.t44 46.4362
R7933 por.n1 por.t30 46.4362
R7934 por.n7 por.t5 39.6005
R7935 por.n7 por.t14 39.6005
R7936 por.n11 por.t7 39.6005
R7937 por.n11 por.t3 39.6005
R7938 por.n15 por.t11 39.6005
R7939 por.n15 por.t15 39.6005
R7940 por.n19 por.t8 39.6005
R7941 por.n19 por.t2 39.6005
R7942 por.n23 por.t12 39.6005
R7943 por.n23 por.t6 39.6005
R7944 por.n27 por.t0 39.6005
R7945 por.n27 por.t9 39.6005
R7946 por.n31 por.t4 39.6005
R7947 por.n31 por.t13 39.6005
R7948 por.n3 por.t1 39.6005
R7949 por.n3 por.t10 39.6005
R7950 por.n40 por 2.2419
R7951 por.n38 por.n6 0.504406
R7952 por.n37 por.n10 0.504406
R7953 por.n36 por.n14 0.504406
R7954 por.n35 por.n18 0.504406
R7955 por.n34 por.n22 0.504406
R7956 por.n33 por.n26 0.504406
R7957 por.n32 por.n30 0.504406
R7958 por.n39 por.n2 0.494641
R7959 por.n38 por.n37 0.276362
R7960 por.n37 por.n36 0.276362
R7961 por.n36 por.n35 0.276362
R7962 por.n35 por.n34 0.276362
R7963 por.n34 por.n33 0.276362
R7964 por.n33 por.n32 0.276362
R7965 por.n39 por.n38 0.267768
R7966 por por.n39 0.187416
R7967 por.n40 por 0.121995
R7968 por por.n40 0.06425
R7969 x2.vbp1.n8 x2.vbp1.t29 231.19
R7970 x2.vbp1.n8 x2.vbp1.t28 230.76
R7971 x2.vbp1.n12 x2.vbp1.n11 202.703
R7972 x2.vbp1.n0 x2.vbp1.n9 202.363
R7973 x2.vbp1.n12 x2.vbp1.n10 202.169
R7974 x2.vbp1.n0 x2.vbp1.n13 201.992
R7975 x2.vbp1.n15 x2.vbp1.n14 201.984
R7976 x2.vbp1.n17 x2.vbp1.n16 201.984
R7977 x2.vbp1.n19 x2.vbp1.n18 201.984
R7978 x2.vbp1.n31 x2.vbp1.t26 121.873
R7979 x2.vbp1.n4 x2.vbp1.t18 121.773
R7980 x2.vbp1.n3 x2.vbp1.t10 121.773
R7981 x2.vbp1.n2 x2.vbp1.t8 121.773
R7982 x2.vbp1.n26 x2.vbp1.t14 121.773
R7983 x2.vbp1.n27 x2.vbp1.t20 121.773
R7984 x2.vbp1.n28 x2.vbp1.t4 121.773
R7985 x2.vbp1.n29 x2.vbp1.t24 121.773
R7986 x2.vbp1.n30 x2.vbp1.t16 121.773
R7987 x2.vbp1.n6 x2.vbp1.t6 121.773
R7988 x2.vbp1.n5 x2.vbp1.t12 121.773
R7989 x2.vbp1.n7 x2.vbp1.t39 121.38
R7990 x2.vbp1.n31 x2.vbp1.t0 121.24
R7991 x2.vbp1.n7 x2.vbp1.t31 120.772
R7992 x2.vbp1.n4 x2.vbp1.t32 119.876
R7993 x2.vbp1.n3 x2.vbp1.t35 119.876
R7994 x2.vbp1.n2 x2.vbp1.t36 119.876
R7995 x2.vbp1.n26 x2.vbp1.t33 119.876
R7996 x2.vbp1.n27 x2.vbp1.t40 119.876
R7997 x2.vbp1.n28 x2.vbp1.t38 119.876
R7998 x2.vbp1.n29 x2.vbp1.t2 119.876
R7999 x2.vbp1.n30 x2.vbp1.t22 119.876
R8000 x2.vbp1.n6 x2.vbp1.t37 119.876
R8001 x2.vbp1.n5 x2.vbp1.t34 119.876
R8002 x2.vbp1.n9 x2.vbp1.t25 28.5655
R8003 x2.vbp1.n9 x2.vbp1.t17 28.5655
R8004 x2.vbp1.n13 x2.vbp1.t21 28.5655
R8005 x2.vbp1.n13 x2.vbp1.t5 28.5655
R8006 x2.vbp1.n14 x2.vbp1.t9 28.5655
R8007 x2.vbp1.n14 x2.vbp1.t15 28.5655
R8008 x2.vbp1.n16 x2.vbp1.t19 28.5655
R8009 x2.vbp1.n16 x2.vbp1.t11 28.5655
R8010 x2.vbp1.n18 x2.vbp1.t7 28.5655
R8011 x2.vbp1.n18 x2.vbp1.t13 28.5655
R8012 x2.vbp1.n10 x2.vbp1.t3 28.5655
R8013 x2.vbp1.n10 x2.vbp1.t23 28.5655
R8014 x2.vbp1.n11 x2.vbp1.t1 28.5655
R8015 x2.vbp1.n11 x2.vbp1.t27 28.5655
R8016 x2.vbp1.n1 x2.vbp1.t30 20.641
R8017 x2.vbp1.n0 x2.vbp1.n12 10.2798
R8018 x2.vbp1.n1 x2.vbp1.n21 3.14057
R8019 x2.vbp1.n32 x2.vbp1.n31 1.56905
R8020 x2.vbp1.n25 x2.vbp1.n24 1.56502
R8021 x2.vbp1.n23 x2.vbp1.n22 1.56194
R8022 x2.vbp1.n34 x2.vbp1.n33 1.54889
R8023 x2.vbp1 x2.vbp1.n35 1.53679
R8024 x2.vbp1.n23 x2.vbp1.n4 1.36443
R8025 x2.vbp1.n24 x2.vbp1.n3 1.36443
R8026 x2.vbp1.n25 x2.vbp1.n2 1.36443
R8027 x2.vbp1 x2.vbp1.n26 1.36443
R8028 x2.vbp1.n35 x2.vbp1.n27 1.36443
R8029 x2.vbp1.n34 x2.vbp1.n28 1.36443
R8030 x2.vbp1.n33 x2.vbp1.n29 1.36443
R8031 x2.vbp1.n32 x2.vbp1.n30 1.36443
R8032 x2.vbp1.n1 x2.vbp1.n6 1.3362
R8033 x2.vbp1.n22 x2.vbp1.n5 1.3362
R8034 x2.vbp1.n21 x2.vbp1.n20 1.33294
R8035 x2.vbp1.n15 x2.vbp1.n0 1.04868
R8036 x2.vbp1.n19 x2.vbp1.n17 0.707531
R8037 x2.vbp1.n17 x2.vbp1.n15 0.707531
R8038 x2.vbp1.n21 x2.vbp1.n7 0.690016
R8039 x2.vbp1.n35 x2.vbp1.n34 0.657758
R8040 x2.vbp1.n33 x2.vbp1.n32 0.641629
R8041 x2.vbp1.n24 x2.vbp1.n23 0.637597
R8042 x2.vbp1 x2.vbp1.n25 0.637597
R8043 x2.vbp1.n20 x2.vbp1.n8 0.601259
R8044 x2.vbp1.n22 x2.vbp1.n1 0.493921
R8045 x2.vbp1.n20 x2.vbp1.n19 0.493624
R8046 a_28094_n290278.n1 a_28094_n290278.t9 231.464
R8047 a_28094_n290278.n1 a_28094_n290278.t8 230.524
R8048 a_28094_n290278.n5 a_28094_n290278.n4 202.834
R8049 a_28094_n290278.n2 a_28094_n290278.n0 202.144
R8050 a_28094_n290278.n7 a_28094_n290278.n6 202.126
R8051 a_28094_n290278.n5 a_28094_n290278.n3 202.112
R8052 a_28094_n290278.n4 a_28094_n290278.t0 28.5655
R8053 a_28094_n290278.n4 a_28094_n290278.t1 28.5655
R8054 a_28094_n290278.n0 a_28094_n290278.t2 28.5655
R8055 a_28094_n290278.n0 a_28094_n290278.t5 28.5655
R8056 a_28094_n290278.n3 a_28094_n290278.t3 28.5655
R8057 a_28094_n290278.n3 a_28094_n290278.t6 28.5655
R8058 a_28094_n290278.t7 a_28094_n290278.n7 28.5655
R8059 a_28094_n290278.n7 a_28094_n290278.t4 28.5655
R8060 a_28094_n290278.n2 a_28094_n290278.n1 1.35637
R8061 a_28094_n290278.n6 a_28094_n290278.n2 0.703306
R8062 a_28094_n290278.n6 a_28094_n290278.n5 0.673969
R8063 x1.vt x1.vt.t3 196.327
R8064 x1.vt.n0 x1.vt.t2 61.721
R8065 x1.vt.n0 x1.vt.t0 25.6927
R8066 x1.vt x1.vt.t1 3.36884
R8067 x1.vt x1.vt.n0 2.46171
R8068 x1.vo.n0 x1.vo.t4 191.04
R8069 x1.vo.n0 x1.vo.t3 123.525
R8070 x1.vo.n3 x1.vo.t2 62.0831
R8071 x1.vo.n2 x1.vo.t1 42.0629
R8072 x1.vo.n2 x1.vo.t0 40.9588
R8073 x1.vo.n1 x1.vo.t5 3.04868
R8074 x1.vo.n1 x1.vo.n0 1.69203
R8075 x1.vo.n3 x1.vo.n1 1.33861
R8076 x1.vo.n3 x1.vo.n2 1.16907
R8077 a_35469_n289052.t60 a_35469_n289052.t37 353.467
R8078 a_35469_n289052.t39 a_35469_n289052.t64 353.467
R8079 a_35469_n289052.t67 a_35469_n289052.t44 353.467
R8080 a_35469_n289052.t30 a_35469_n289052.t55 353.467
R8081 a_35469_n289052.t56 a_35469_n289052.t36 353.467
R8082 a_35469_n289052.t41 a_35469_n289052.t69 353.467
R8083 a_35469_n289052.t70 a_35469_n289052.t46 353.467
R8084 a_35469_n289052.t48 a_35469_n289052.t26 353.467
R8085 a_35469_n289052.t35 a_35469_n289052.t58 353.467
R8086 a_35469_n289052.t40 a_35469_n289052.t68 353.467
R8087 a_35469_n289052.t25 a_35469_n289052.t50 353.467
R8088 a_35469_n289052.t52 a_35469_n289052.t31 353.467
R8089 a_35469_n289052.t33 a_35469_n289052.t57 353.467
R8090 a_35469_n289052.t65 a_35469_n289052.t42 353.467
R8091 a_35469_n289052.t45 a_35469_n289052.t71 353.467
R8092 a_35469_n289052.t29 a_35469_n289052.t53 353.467
R8093 a_35469_n289052.n0 a_35469_n289052.n10 299.851
R8094 a_35469_n289052.n0 a_35469_n289052.n7 299.851
R8095 a_35469_n289052.n1 a_35469_n289052.n4 299.851
R8096 a_35469_n289052.n44 a_35469_n289052.n1 299.851
R8097 a_35469_n289052.n1 a_35469_n289052.n43 299.414
R8098 a_35469_n289052.n0 a_35469_n289052.n11 299.414
R8099 a_35469_n289052.n0 a_35469_n289052.n8 299.414
R8100 a_35469_n289052.n1 a_35469_n289052.n5 299.414
R8101 a_35469_n289052.n34 a_35469_n289052.t60 232.382
R8102 a_35469_n289052.n27 a_35469_n289052.t29 232.382
R8103 a_35469_n289052.n1 a_35469_n289052.n2 197.123
R8104 a_35469_n289052.n0 a_35469_n289052.n9 197.123
R8105 a_35469_n289052.n0 a_35469_n289052.n6 197.123
R8106 a_35469_n289052.n1 a_35469_n289052.n3 197.123
R8107 a_35469_n289052.n12 a_35469_n289052.t49 185.79
R8108 a_35469_n289052.n19 a_35469_n289052.t34 185.79
R8109 a_35469_n289052.n34 a_35469_n289052.t39 162.274
R8110 a_35469_n289052.n35 a_35469_n289052.t67 162.274
R8111 a_35469_n289052.n36 a_35469_n289052.t30 162.274
R8112 a_35469_n289052.n37 a_35469_n289052.t56 162.274
R8113 a_35469_n289052.n38 a_35469_n289052.t41 162.274
R8114 a_35469_n289052.n39 a_35469_n289052.t70 162.274
R8115 a_35469_n289052.n40 a_35469_n289052.t48 162.274
R8116 a_35469_n289052.n33 a_35469_n289052.t35 162.274
R8117 a_35469_n289052.n32 a_35469_n289052.t40 162.274
R8118 a_35469_n289052.n31 a_35469_n289052.t25 162.274
R8119 a_35469_n289052.n30 a_35469_n289052.t52 162.274
R8120 a_35469_n289052.n29 a_35469_n289052.t33 162.274
R8121 a_35469_n289052.n28 a_35469_n289052.t65 162.274
R8122 a_35469_n289052.n27 a_35469_n289052.t45 162.274
R8123 a_35469_n289052.n12 a_35469_n289052.t66 115.68
R8124 a_35469_n289052.n13 a_35469_n289052.t38 115.68
R8125 a_35469_n289052.n14 a_35469_n289052.t59 115.68
R8126 a_35469_n289052.n15 a_35469_n289052.t27 115.68
R8127 a_35469_n289052.n16 a_35469_n289052.t47 115.68
R8128 a_35469_n289052.n17 a_35469_n289052.t62 115.68
R8129 a_35469_n289052.n18 a_35469_n289052.t54 115.68
R8130 a_35469_n289052.n25 a_35469_n289052.t28 115.68
R8131 a_35469_n289052.n24 a_35469_n289052.t43 115.68
R8132 a_35469_n289052.n23 a_35469_n289052.t63 115.68
R8133 a_35469_n289052.n22 a_35469_n289052.t32 115.68
R8134 a_35469_n289052.n21 a_35469_n289052.t51 115.68
R8135 a_35469_n289052.n20 a_35469_n289052.t24 115.68
R8136 a_35469_n289052.n19 a_35469_n289052.t61 115.68
R8137 a_35469_n289052.n28 a_35469_n289052.n27 70.1096
R8138 a_35469_n289052.n29 a_35469_n289052.n28 70.1096
R8139 a_35469_n289052.n30 a_35469_n289052.n29 70.1096
R8140 a_35469_n289052.n31 a_35469_n289052.n30 70.1096
R8141 a_35469_n289052.n32 a_35469_n289052.n31 70.1096
R8142 a_35469_n289052.n33 a_35469_n289052.n32 70.1096
R8143 a_35469_n289052.n40 a_35469_n289052.n39 70.1096
R8144 a_35469_n289052.n39 a_35469_n289052.n38 70.1096
R8145 a_35469_n289052.n38 a_35469_n289052.n37 70.1096
R8146 a_35469_n289052.n37 a_35469_n289052.n36 70.1096
R8147 a_35469_n289052.n36 a_35469_n289052.n35 70.1096
R8148 a_35469_n289052.n35 a_35469_n289052.n34 70.1096
R8149 a_35469_n289052.n13 a_35469_n289052.n12 70.1096
R8150 a_35469_n289052.n14 a_35469_n289052.n13 70.1096
R8151 a_35469_n289052.n15 a_35469_n289052.n14 70.1096
R8152 a_35469_n289052.n16 a_35469_n289052.n15 70.1096
R8153 a_35469_n289052.n17 a_35469_n289052.n16 70.1096
R8154 a_35469_n289052.n18 a_35469_n289052.n17 70.1096
R8155 a_35469_n289052.n25 a_35469_n289052.n24 70.1096
R8156 a_35469_n289052.n24 a_35469_n289052.n23 70.1096
R8157 a_35469_n289052.n23 a_35469_n289052.n22 70.1096
R8158 a_35469_n289052.n22 a_35469_n289052.n21 70.1096
R8159 a_35469_n289052.n21 a_35469_n289052.n20 70.1096
R8160 a_35469_n289052.n20 a_35469_n289052.n19 70.1096
R8161 a_35469_n289052.n43 a_35469_n289052.t6 46.4362
R8162 a_35469_n289052.n43 a_35469_n289052.t2 46.4362
R8163 a_35469_n289052.n11 a_35469_n289052.t21 46.4362
R8164 a_35469_n289052.n11 a_35469_n289052.t12 46.4362
R8165 a_35469_n289052.n10 a_35469_n289052.t17 46.4362
R8166 a_35469_n289052.n10 a_35469_n289052.t20 46.4362
R8167 a_35469_n289052.n8 a_35469_n289052.t22 46.4362
R8168 a_35469_n289052.n8 a_35469_n289052.t19 46.4362
R8169 a_35469_n289052.n7 a_35469_n289052.t4 46.4362
R8170 a_35469_n289052.n7 a_35469_n289052.t3 46.4362
R8171 a_35469_n289052.n5 a_35469_n289052.t8 46.4362
R8172 a_35469_n289052.n5 a_35469_n289052.t1 46.4362
R8173 a_35469_n289052.n4 a_35469_n289052.t18 46.4362
R8174 a_35469_n289052.n4 a_35469_n289052.t10 46.4362
R8175 a_35469_n289052.t0 a_35469_n289052.n44 46.4362
R8176 a_35469_n289052.n44 a_35469_n289052.t14 46.4362
R8177 a_35469_n289052.n2 a_35469_n289052.t23 39.6005
R8178 a_35469_n289052.n2 a_35469_n289052.t15 39.6005
R8179 a_35469_n289052.n9 a_35469_n289052.t13 39.6005
R8180 a_35469_n289052.n9 a_35469_n289052.t11 39.6005
R8181 a_35469_n289052.n6 a_35469_n289052.t5 39.6005
R8182 a_35469_n289052.n6 a_35469_n289052.t9 39.6005
R8183 a_35469_n289052.n3 a_35469_n289052.t16 39.6005
R8184 a_35469_n289052.n3 a_35469_n289052.t7 39.6005
R8185 a_35469_n289052.n41 a_35469_n289052.n33 35.055
R8186 a_35469_n289052.n41 a_35469_n289052.n40 35.055
R8187 a_35469_n289052.n26 a_35469_n289052.n18 35.055
R8188 a_35469_n289052.n26 a_35469_n289052.n25 35.055
R8189 a_35469_n289052.n42 a_35469_n289052.n26 10.2069
R8190 a_35469_n289052.n42 a_35469_n289052.n41 10.156
R8191 a_35469_n289052.n1 a_35469_n289052.n0 2.84371
R8192 a_35469_n289052.n0 a_35469_n289052.n42 2.6231
R8193 porb.n7 porb.n5 299.851
R8194 porb.n11 porb.n9 299.851
R8195 porb.n15 porb.n13 299.851
R8196 porb.n19 porb.n17 299.851
R8197 porb.n23 porb.n21 299.851
R8198 porb.n27 porb.n25 299.851
R8199 porb.n31 porb.n29 299.851
R8200 porb.n3 porb.n1 299.851
R8201 porb.n7 porb.n6 299.414
R8202 porb.n11 porb.n10 299.414
R8203 porb.n15 porb.n14 299.414
R8204 porb.n19 porb.n18 299.414
R8205 porb.n23 porb.n22 299.414
R8206 porb.n27 porb.n26 299.414
R8207 porb.n31 porb.n30 299.414
R8208 porb.n3 porb.n2 299.414
R8209 porb.n38 porb.n4 197.123
R8210 porb.n37 porb.n8 197.123
R8211 porb.n36 porb.n12 197.123
R8212 porb.n35 porb.n16 197.123
R8213 porb.n34 porb.n20 197.123
R8214 porb.n33 porb.n24 197.123
R8215 porb.n32 porb.n28 197.123
R8216 porb.n39 porb.n0 197.094
R8217 porb.n6 porb.t21 46.4362
R8218 porb.n6 porb.t42 46.4362
R8219 porb.n5 porb.t35 46.4362
R8220 porb.n5 porb.t25 46.4362
R8221 porb.n10 porb.t29 46.4362
R8222 porb.n10 porb.t47 46.4362
R8223 porb.n9 porb.t43 46.4362
R8224 porb.n9 porb.t30 46.4362
R8225 porb.n14 porb.t37 46.4362
R8226 porb.n14 porb.t41 46.4362
R8227 porb.n13 porb.t19 46.4362
R8228 porb.n13 porb.t24 46.4362
R8229 porb.n18 porb.t31 46.4362
R8230 porb.n18 porb.t17 46.4362
R8231 porb.n17 porb.t46 46.4362
R8232 porb.n17 porb.t32 46.4362
R8233 porb.n22 porb.t36 46.4362
R8234 porb.n22 porb.t26 46.4362
R8235 porb.n21 porb.t18 46.4362
R8236 porb.n21 porb.t40 46.4362
R8237 porb.n26 porb.t44 46.4362
R8238 porb.n26 porb.t20 46.4362
R8239 porb.n25 porb.t27 46.4362
R8240 porb.n25 porb.t34 46.4362
R8241 porb.n30 porb.t38 46.4362
R8242 porb.n30 porb.t23 46.4362
R8243 porb.n29 porb.t22 46.4362
R8244 porb.n29 porb.t39 46.4362
R8245 porb.n2 porb.t45 46.4362
R8246 porb.n2 porb.t33 46.4362
R8247 porb.n1 porb.t28 46.4362
R8248 porb.n1 porb.t16 46.4362
R8249 porb.n4 porb.t10 39.6005
R8250 porb.n4 porb.t4 39.6005
R8251 porb.n8 porb.t14 39.6005
R8252 porb.n8 porb.t8 39.6005
R8253 porb.n12 porb.t2 39.6005
R8254 porb.n12 porb.t5 39.6005
R8255 porb.n16 porb.t13 39.6005
R8256 porb.n16 porb.t9 39.6005
R8257 porb.n20 porb.t1 39.6005
R8258 porb.n20 porb.t12 39.6005
R8259 porb.n24 porb.t6 39.6005
R8260 porb.n24 porb.t15 39.6005
R8261 porb.n28 porb.t3 39.6005
R8262 porb.n28 porb.t11 39.6005
R8263 porb.n0 porb.t7 39.6005
R8264 porb.n0 porb.t0 39.6005
R8265 porb.n38 porb.n7 0.504406
R8266 porb.n37 porb.n11 0.504406
R8267 porb.n36 porb.n15 0.504406
R8268 porb.n35 porb.n19 0.504406
R8269 porb.n34 porb.n23 0.504406
R8270 porb.n33 porb.n27 0.504406
R8271 porb.n32 porb.n31 0.504406
R8272 porb.n39 porb.n3 0.494641
R8273 porb.n38 porb.n37 0.276362
R8274 porb.n37 porb.n36 0.276362
R8275 porb.n36 porb.n35 0.276362
R8276 porb.n35 porb.n34 0.276362
R8277 porb.n34 porb.n33 0.276362
R8278 porb.n33 porb.n32 0.276362
R8279 porb.n39 porb.n38 0.267768
R8280 porb porb.n39 0.254005
R8281 a_35277_n289052.t10 a_35277_n289052.t22 353.467
R8282 a_35277_n289052.t26 a_35277_n289052.t14 353.467
R8283 a_35277_n289052.t15 a_35277_n289052.t28 353.467
R8284 a_35277_n289052.t8 a_35277_n289052.t20 353.467
R8285 a_35277_n289052.t21 a_35277_n289052.t11 353.467
R8286 a_35277_n289052.t12 a_35277_n289052.t24 353.467
R8287 a_35277_n289052.t16 a_35277_n289052.t6 353.467
R8288 a_35277_n289052.t7 a_35277_n289052.t19 353.467
R8289 a_35277_n289052.n18 a_35277_n289052.n17 299.851
R8290 a_35277_n289052.n19 a_35277_n289052.n18 299.414
R8291 a_35277_n289052.n11 a_35277_n289052.t10 232.382
R8292 a_35277_n289052.n8 a_35277_n289052.t7 232.382
R8293 a_35277_n289052.n16 a_35277_n289052.n0 197.161
R8294 a_35277_n289052.n1 a_35277_n289052.t17 185.79
R8295 a_35277_n289052.n4 a_35277_n289052.t23 185.79
R8296 a_35277_n289052.n11 a_35277_n289052.t26 162.274
R8297 a_35277_n289052.n12 a_35277_n289052.t15 162.274
R8298 a_35277_n289052.n13 a_35277_n289052.t8 162.274
R8299 a_35277_n289052.n10 a_35277_n289052.t21 162.274
R8300 a_35277_n289052.n9 a_35277_n289052.t12 162.274
R8301 a_35277_n289052.n8 a_35277_n289052.t16 162.274
R8302 a_35277_n289052.n1 a_35277_n289052.t29 115.68
R8303 a_35277_n289052.n2 a_35277_n289052.t25 115.68
R8304 a_35277_n289052.n3 a_35277_n289052.t9 115.68
R8305 a_35277_n289052.n6 a_35277_n289052.t18 115.68
R8306 a_35277_n289052.n5 a_35277_n289052.t27 115.68
R8307 a_35277_n289052.n4 a_35277_n289052.t13 115.68
R8308 a_35277_n289052.n9 a_35277_n289052.n8 70.1096
R8309 a_35277_n289052.n10 a_35277_n289052.n9 70.1096
R8310 a_35277_n289052.n13 a_35277_n289052.n12 70.1096
R8311 a_35277_n289052.n12 a_35277_n289052.n11 70.1096
R8312 a_35277_n289052.n2 a_35277_n289052.n1 70.1096
R8313 a_35277_n289052.n3 a_35277_n289052.n2 70.1096
R8314 a_35277_n289052.n6 a_35277_n289052.n5 70.1096
R8315 a_35277_n289052.n5 a_35277_n289052.n4 70.1096
R8316 a_35277_n289052.n17 a_35277_n289052.t4 46.4362
R8317 a_35277_n289052.n17 a_35277_n289052.t3 46.4362
R8318 a_35277_n289052.n19 a_35277_n289052.t2 46.4362
R8319 a_35277_n289052.t5 a_35277_n289052.n19 46.4362
R8320 a_35277_n289052.n0 a_35277_n289052.t1 39.6005
R8321 a_35277_n289052.n0 a_35277_n289052.t0 39.6005
R8322 a_35277_n289052.n14 a_35277_n289052.n10 35.055
R8323 a_35277_n289052.n14 a_35277_n289052.n13 35.055
R8324 a_35277_n289052.n7 a_35277_n289052.n3 35.055
R8325 a_35277_n289052.n7 a_35277_n289052.n6 35.055
R8326 a_35277_n289052.n15 a_35277_n289052.n7 17.6874
R8327 a_35277_n289052.n15 a_35277_n289052.n14 17.6491
R8328 a_35277_n289052.n16 a_35277_n289052.n15 2.43319
R8329 a_35277_n289052.n18 a_35277_n289052.n16 0.572285
R8330 x1.Vinn.n3 x1.Vinn.t5 71.5611
R8331 x1.Vinn.n0 x1.Vinn.t2 71.5515
R8332 x1.Vinn.n1 x1.Vinn.t3 71.5483
R8333 x1.Vinn.n3 x1.Vinn.t4 71.3939
R8334 x1.Vinn.n0 x1.Vinn.t6 71.3938
R8335 x1.Vinn.n1 x1.Vinn.t7 71.3918
R8336 x1.Vinn.n5 x1.Vinn.t1 42.6627
R8337 x1.Vinn x1.Vinn.n5 4.7372
R8338 x1.Vinn.n5 x1.Vinn.t0 3.13485
R8339 x1.Vinn.n2 x1.Vinn.n0 2.10424
R8340 x1.Vinn.n2 x1.Vinn.n1 1.1401
R8341 x1.Vinn.n4 x1.Vinn.n3 1.12922
R8342 x1.Vinn.n4 x1.Vinn.n2 1.01093
R8343 x1.Vinn x1.Vinn.n4 0.688261
R8344 a_24270_n290121.n0 a_24270_n290121.t1 114.763
R8345 a_24270_n290121.n4 a_24270_n290121.n2 102.094
R8346 a_24270_n290121.n14 a_24270_n290121.n13 101.809
R8347 a_24270_n290121.n4 a_24270_n290121.n3 101.799
R8348 a_24270_n290121.n12 a_24270_n290121.n11 101.793
R8349 a_24270_n290121.n1 a_24270_n290121.t4 81.3863
R8350 a_24270_n290121.n1 a_24270_n290121.t18 80.9347
R8351 a_24270_n290121.n1 a_24270_n290121.t14 80.6566
R8352 a_24270_n290121.n5 a_24270_n290121.t8 80.6566
R8353 a_24270_n290121.n6 a_24270_n290121.t16 80.6566
R8354 a_24270_n290121.n7 a_24270_n290121.t2 80.6566
R8355 a_24270_n290121.n8 a_24270_n290121.t12 80.6566
R8356 a_24270_n290121.n9 a_24270_n290121.t10 80.6566
R8357 a_24270_n290121.n10 a_24270_n290121.t6 80.6566
R8358 a_24270_n290121.n11 a_24270_n290121.t11 13.848
R8359 a_24270_n290121.n11 a_24270_n290121.t7 13.848
R8360 a_24270_n290121.n3 a_24270_n290121.t9 13.848
R8361 a_24270_n290121.n3 a_24270_n290121.t17 13.848
R8362 a_24270_n290121.n2 a_24270_n290121.t5 13.848
R8363 a_24270_n290121.n2 a_24270_n290121.t15 13.848
R8364 a_24270_n290121.n14 a_24270_n290121.t3 13.848
R8365 a_24270_n290121.t13 a_24270_n290121.n14 13.848
R8366 a_24270_n290121.n0 a_24270_n290121.t0 6.39288
R8367 a_24270_n290121.n0 a_24270_n290121.n10 1.55432
R8368 a_24270_n290121.n6 a_24270_n290121.n5 0.7505
R8369 a_24270_n290121.n9 a_24270_n290121.n8 0.740365
R8370 a_24270_n290121.n7 a_24270_n290121.n6 0.736986
R8371 a_24270_n290121.n10 a_24270_n290121.n9 0.736986
R8372 a_24270_n290121.n8 a_24270_n290121.n7 0.726851
R8373 a_24270_n290121.n5 a_24270_n290121.n1 0.726851
R8374 a_24270_n290121.n12 a_24270_n290121.n0 0.528774
R8375 a_24270_n290121.n13 a_24270_n290121.n12 0.325649
R8376 a_24270_n290121.n13 a_24270_n290121.n4 0.324161
R8377 a_34015_n286994.n3 a_34015_n286994.t4 332.315
R8378 a_34015_n286994.t4 a_34015_n286994.n2 332.296
R8379 a_34015_n286994.n3 a_34015_n286994.t5 331.928
R8380 a_34015_n286994.t5 a_34015_n286994.n2 331.928
R8381 a_34015_n286994.n0 a_34015_n286994.t2 85.8522
R8382 a_34015_n286994.t3 a_34015_n286994.n1 84.1877
R8383 a_34015_n286994.n0 a_34015_n286994.t0 49.8239
R8384 a_34015_n286994.n0 a_34015_n286994.t1 49.8155
R8385 a_34015_n286994.n1 a_34015_n286994.n0 2.13415
R8386 a_34015_n286994.n1 a_34015_n286994.n2 1.74288
R8387 a_34015_n286994.n1 a_34015_n286994.n3 1.15456
R8388 x2.vbn1.n6 x2.vbn1.t15 115.534
R8389 x2.vbn1.n2 x2.vbn1.t16 80.1876
R8390 x2.vbn1.n7 x2.vbn1.t13 79.4015
R8391 x2.vbn1.n8 x2.vbn1.t3 79.4015
R8392 x2.vbn1.n9 x2.vbn1.t5 79.4015
R8393 x2.vbn1.n10 x2.vbn1.t11 79.4015
R8394 x2.vbn1.n11 x2.vbn1.t9 79.4015
R8395 x2.vbn1.n12 x2.vbn1.t1 79.4015
R8396 x2.vbn1.n13 x2.vbn1.t7 79.4015
R8397 x2.vbn1.n14 x2.vbn1.t18 79.4015
R8398 x2.vbn1.n15 x2.vbn1.t17 79.4015
R8399 x2.vbn1.n16 x2.vbn1.t20 79.4015
R8400 x2.vbn1.n2 x2.vbn1.t19 79.4015
R8401 x2.vbn1.n1 x2.vbn1.t14 43.482
R8402 x2.vbn1.n0 x2.vbn1.n3 35.5796
R8403 x2.vbn1.n0 x2.vbn1.n5 35.2408
R8404 x2.vbn1.n0 x2.vbn1.n4 35.2326
R8405 x2.vbn1.n5 x2.vbn1.t6 8.2655
R8406 x2.vbn1.n5 x2.vbn1.t4 8.2655
R8407 x2.vbn1.n4 x2.vbn1.t10 8.2655
R8408 x2.vbn1.n4 x2.vbn1.t12 8.2655
R8409 x2.vbn1.n3 x2.vbn1.t8 8.2655
R8410 x2.vbn1.n3 x2.vbn1.t2 8.2655
R8411 x2.vbn1.n6 x2.vbn1.t0 4.44838
R8412 x2.vbn1.n15 x2.vbn1.n14 1.83506
R8413 x2.vbn1.n14 x2.vbn1.n13 1.80197
R8414 x2.vbn1.n7 x2.vbn1.n1 1.67073
R8415 x2.vbn1.n1 x2.vbn1.n6 1.18037
R8416 x2.vbn1.n1 x2.vbn1.n0 0.867602
R8417 x2.vbn1.n16 x2.vbn1.n15 0.827706
R8418 x2.vbn1.n13 x2.vbn1.n12 0.813
R8419 x2.vbn1.n12 x2.vbn1.n11 0.809324
R8420 x2.vbn1.n10 x2.vbn1.n9 0.809324
R8421 x2.vbn1.n8 x2.vbn1.n7 0.805647
R8422 x2.vbn1.n9 x2.vbn1.n8 0.794618
R8423 x2.vbn1.n11 x2.vbn1.n10 0.787265
R8424 x2.vbn1.n16 x2.vbn1.n2 0.776235
R8425 a_13449_n292106.n0 a_13449_n292106.t3 194.236
R8426 a_13449_n292106.n0 a_13449_n292106.t1 193.607
R8427 a_13449_n292106.t2 a_13449_n292106.n0 61.7906
R8428 a_13449_n292106.n0 a_13449_n292106.t0 25.6009
R8429 x2.x3.aout.n1 x2.x3.aout.t3 157.346
R8430 x2.x3.aout.n1 x2.x3.aout.t4 157.346
R8431 x2.x3.aout.n1 x2.x3.aout.t5 119.2
R8432 x2.x3.aout.n1 x2.x3.aout.t6 119.2
R8433 x2.x3.aout.n0 x2.x3.aout.t1 85.7689
R8434 x2.x3.aout.n0 x2.x3.aout.t2 85.6122
R8435 x2.x3.aout.n0 x2.x3.aout.t0 49.7738
R8436 x2.x3.aout.n0 x2.x3.aout 12.5005
R8437 x2.x3.aout.n0 x2.x3.aout.n1 2.97733
R8438 x1.VD.n2 x1.VD.t0 113.207
R8439 x1.VD.n2 x1.VD.t2 84.8264
R8440 x1.VD.n1 x1.VD.t8 43.9926
R8441 x1.VD.n0 x1.VD.t7 43.9576
R8442 x1.VD.n1 x1.VD.t3 43.8803
R8443 x1.VD.n1 x1.VD.t6 43.8696
R8444 x1.VD.n0 x1.VD.t4 43.856
R8445 x1.VD.n0 x1.VD.t5 43.8457
R8446 x1.VD x1.VD.t1 23.5777
R8447 x1.VD.n4 x1.VD.n0 3.71432
R8448 x1.VD x1.VD.n4 3.45953
R8449 x1.VD.n3 x1.VD 3.28686
R8450 x1.VD.n3 x1.VD.n0 3.03806
R8451 x1.VD.n4 x1.VD.n1 3.02208
R8452 x1.VD.n1 x1.VD.n3 2.35302
R8453 x1.VD x1.VD.n2 1.60343
R8454 a_24253_n287224.n1 a_24253_n287224.t10 145.53
R8455 a_24253_n287224.n1 a_24253_n287224.n3 2.12261
R8456 a_24253_n287224.t9 a_24253_n287224.n3 128.244
R8457 a_24253_n287224.n0 a_24253_n287224.t4 128.24
R8458 a_24253_n287224.t6 a_24253_n287224.n3 128.048
R8459 a_24253_n287224.t11 a_24253_n287224.n0 128.048
R8460 a_24253_n287224.n5 a_24253_n287224.n0 5.60863
R8461 a_24253_n287224.n2 a_24253_n287224.t0 232.814
R8462 a_24253_n287224.n2 a_24253_n287224.t1 232.075
R8463 a_24253_n287224.n1 a_24253_n287224.t2 228.215
R8464 a_24253_n287224.t3 a_24253_n287224.n1 228.215
R8465 a_24253_n287224.n1 a_24253_n287224.t8 146.207
R8466 a_24253_n287224.n4 a_24253_n287224.t7 145.499
R8467 a_24253_n287224.n4 a_24253_n287224.t5 145.316
R8468 a_24253_n287224.n1 a_24253_n287224.n5 28.2118
R8469 a_24253_n287224.n5 a_24253_n287224.n4 3.66328
R8470 a_24253_n287224.n1 a_24253_n287224.n2 3.42195
R8471 x2.Td_S x2.Td_S.t1 232.379
R8472 x2.Td_S x2.Td_S.t0 232.141
R8473 x2.Td_S x2.Td_S.t3 231.448
R8474 x2.Td_S x2.Td_S.t2 230.472
R8475 x2.Td_S.n0 x2.Td_S.t6 175.066
R8476 x2.Td_S.n0 x2.Td_S.t4 173.9
R8477 x2.Td_S.n0 x2.Td_S.t5 164.5
R8478 x2.Td_S x2.Td_S.n0 4.55127
R8479 a_24570_n290925.t3 a_24570_n290925.n0 113.207
R8480 a_24570_n290925.n1 a_24570_n290925.t1 86.2485
R8481 a_24570_n290925.n0 a_24570_n290925.t4 81.5196
R8482 a_24570_n290925.n0 a_24570_n290925.t2 80.9292
R8483 a_24570_n290925.n0 a_24570_n290925.n1 3.10362
R8484 a_24570_n290925.n1 a_24570_n290925.t0 2.49272
R8485 x1.Vinp.n0 x1.Vinp.t3 71.5399
R8486 x1.Vinp.n0 x1.Vinp.t2 71.3958
R8487 x1.Vinp.n1 x1.Vinp.t1 42.4766
R8488 x1.Vinp.n1 x1.Vinp.t0 42.4696
R8489 x1.Vinp x1.Vinp.n1 11.3625
R8490 x1.Vinp x1.Vinp.n0 6.32021
R8491 a_4508_n291419.t0 a_4508_n291419.t2 228.155
R8492 a_4508_n291419.t1 a_4508_n291419.t0 227.583
R8493 a_4566_n290308.t1 a_4566_n290308.t0 228.111
R8494 a_4566_n290308.t2 a_4566_n290308.t1 227.607
R8495 x1.vo1.n0 x1.vo1.t1 227.345
R8496 x1.vo1.n2 x1.vo1.t6 150.98
R8497 x1.x1.S x1.vo1.t7 145.46
R8498 x1.vo1.n2 x1.vo1.t2 122.59
R8499 x1.vo1.n0 x1.vo1.t5 121.273
R8500 x1.vo1.n1 x1.vo1.t8 120.938
R8501 x1.vo1.n1 x1.vo1.t4 120.442
R8502 x1.x1.S x1.vo1.t3 119.079
R8503 x1.vo1.n3 x1.vo1.t0 21.7966
R8504 x1.vo1.n3 x1.x1.S 16.6411
R8505 x1.vo1.n0 x1.vo1.n1 5.75907
R8506 x1.x1.S x1.vo1.n2 2.65106
R8507 x1.vo1.n3 x1.vo1.n0 2.01423
R8508 x1.VY x1.VY.t3 114.275
R8509 x1.VY.n0 x1.VY.t0 114.109
R8510 x1.VY x1.VY.t1 83.74
R8511 x1.VY.n0 x1.VY.t2 83.529
R8512 x1.VY.n1 x1.VY.t5 46.9976
R8513 x1.VY x1.VY.t4 44.3856
R8514 x1.VY x1.VY.t6 43.954
R8515 x1.VY x1.VY.n1 8.1227
R8516 x1.VY x1.VY.n0 2.82848
R8517 x1.VY.n1 x1.VY 2.36831
R8518 vbg vbg.t0 60.1284
C0 x2.vbp2 dvdd 1.88695f
C1 avdd a_14970_n288829# 0.338226f
C2 x1.VD a_13030_n290763# 0.175334f
C3 x2.Td_Lb a_29671_n288104# 0.155734f
C4 avss w_15901_n291463# 0.524278f
C5 avdd x2.x3.S1B 0.190118f
C6 x2.VT2 a_29688_n287709# 0.023054f
C7 x2.VT3 avss 0.625952f
C8 a_12978_n288829# x1.vt 0.03595f
C9 a_8104_n286429# a_8436_n286429# 0.307869f
C10 avdd dvdd 16.293201f
C11 avdd a_29487_n288398# 0.029396f
C12 x2.Td_S avdd 1.05661f
C13 a_29671_n288104# a_30011_n288135# 0.240541f
C14 a_30699_n288291# dvdd 0.277431f
C15 a_29487_n288398# a_30699_n288291# 0.077664f
C16 porb_h[0] porb_h[1] 0.134177f
C17 x2.Td_L x2.VT2 0.315185f
C18 a_14472_n286429# a_14804_n286429# 0.308171f
C19 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtp_1_0.D a_29211_n288416# 0.186688f
C20 x1.vbn a_8656_n292108# 0.150633f
C21 x2.din a_23173_n289908# 0.077946f
C22 a_25216_n290828# avdd 0.405546f
C23 a_18492_n288774# a_18960_n288774# 0.309677f
C24 a_22471_n292308# vbg 0.05381f
C25 a_29876_n288037# dvdd 0.277611f
C26 x1.Vinp a_12646_n288829# 0.083378f
C27 a_21534_n286374# a_22002_n286374# 0.307869f
C28 a_29487_n288398# a_29876_n288037# 0.060227f
C29 a_30112_n289746# x2.vbp2 0.37558f
C30 x2.vbp1 a_30814_n289746# 0.012704f
C31 a_29214_n287320# a_29481_n287384# 0.279149f
C32 a_18025_n289908# a_18493_n289908# 0.309071f
C33 a_15914_n289870# dvdd 1.15506f
C34 a_10760_n286429# a_11092_n286429# 0.307869f
C35 a_30112_n289746# avdd 0.533657f
C36 a_22003_n292308# vbg 0.05381f
C37 a_20832_n288774# a_21300_n288774# 0.309677f
C38 avdd x2.Td_Lb 0.977643f
C39 a_18960_n288774# x2.din 0.045459f
C40 x2.Td_Lb a_30699_n288291# 0.173535f
C41 a_9266_n288829# a_9598_n288829# 0.307869f
C42 x1.VD x1.vt 0.207045f
C43 x1.VS x1.VD 3.5535f
C44 avss a_10926_n288829# 0.239853f
C45 a_19662_n286374# avdd 0.110373f
C46 x2.din a_18493_n289908# 0.049162f
C47 x2.din a_19429_n289908# 0.042963f
C48 a_17791_n292308# vbg 0.05381f
C49 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtp_1_0.D a_28056_n288420# 0.235129f
C50 a_19896_n288774# dvdd 0.041197f
C51 x2.VT2 a_29895_n287373# 0.031579f
C52 avss a_8436_n286429# 0.197326f
C53 avdd a_30011_n288135# 0.036572f
C54 a_30814_n289746# dvdd 0.328379f
C55 a_29671_n288104# a_30447_n288420# 0.357796f
C56 avss a_14804_n286429# 0.460997f
C57 a_31045_n288085# dvdd 0.213157f
C58 x2.Td_Lb a_29876_n288037# 0.232063f
C59 x2.VT2 a_10096_n286429# 0.013124f
C60 avss a_13030_n290763# 1.02651f
C61 a_32248_n290278# avdd 0.959785f
C62 a_35074_n291454# dvdd 1.29046f
C63 a_18726_n286374# a_19194_n286374# 0.307869f
C64 avss a_9598_n288829# 0.335767f
C65 a_30011_n288135# a_29876_n288037# 0.356154f
C66 x2.porbPre a_35089_n289052# 0.521153f
C67 a_13310_n288829# a_13642_n288829# 0.310806f
C68 a_20599_n292308# a_21067_n292308# 0.309071f
C69 a_30779_n287655# a_31115_n287366# 0.142416f
C70 a_29481_n287384# a_30447_n287429# 0.137783f
C71 a_29688_n287709# a_30779_n287655# 0.034711f
C72 a_21300_n288774# dvdd 0.041197f
C73 x2.vbp1 porb 0.115435f
C74 x2.Td_L x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N 0.035305f
C75 a_10262_n288829# x1.Vinn 0.021375f
C76 avss a_13642_n288829# 0.335953f
C77 a_30112_n289746# a_30814_n289746# 0.267049f
C78 a_21066_n286374# a_21534_n286374# 0.307869f
C79 a_9432_n286429# a_9764_n286429# 0.307869f
C80 x1.VY x1.VS 1.28069f
C81 avss a_8490_n290308# 0.556388f
C82 avss a_12812_n286429# 0.203435f
C83 a_22704_n288774# avdd 0.013837f
C84 a_13310_n288829# x1.vt 0.088384f
C85 x2.vbp2 a_30410_n291353# 0.139528f
C86 avdd a_30447_n288420# 0.060569f
C87 x2.VT2 a_29671_n288104# 0.014487f
C88 a_30699_n288291# a_30447_n288420# 0.273876f
C89 avdd por 0.199947f
C90 a_20364_n288774# a_20832_n288774# 0.309677f
C91 w_15901_n291463# x1.vt 0.307709f
C92 dvdd porb 11.4196f
C93 avdd x2.x3.aout 3.00683f
C94 avss x1.vt 4.55005f
C95 a_30410_n291353# avdd 0.557082f
C96 avss x1.VS 2.63489f
C97 a_22939_n292308# vbg 0.05381f
C98 a_11424_n286429# x1.Vinp 0.031564f
C99 a_28607_n287397# a_28571_n287754# 0.011144f
C100 a_13476_n286429# a_13808_n286429# 0.310806f
C101 a_20833_n289908# a_21301_n289908# 0.309071f
C102 avss a_10096_n286429# 0.197326f
C103 a_30022_n287538# a_30447_n287429# 0.038205f
C104 a_28607_n287397# dvdd 0.234404f
C105 a_29481_n287384# a_30022_n287538# 0.145305f
C106 a_7996_n292010# a_8656_n292108# 0.32514f
C107 x1.vbn x1.VD 0.048231f
C108 a_29214_n287320# dvdd 0.303686f
C109 x2.porbPre dvdd 1.96253f
C110 x2.vbp2 x2.VT2 0.162666f
C111 a_19428_n288774# x2.din 0.045459f
C112 avdd x1.VD 1.32524f
C113 avss a_11258_n288829# 0.240383f
C114 x2.din a_18961_n289908# 0.042963f
C115 a_20130_n286374# avdd 0.110373f
C116 x2.din a_19897_n289908# 0.042963f
C117 a_20364_n288774# dvdd 0.041197f
C118 a_18259_n292308# vbg 0.05381f
C119 a_19195_n292308# vbg 0.05381f
C120 avss a_8768_n286429# 0.197326f
C121 a_8270_n288829# a_8602_n288829# 0.307869f
C122 x2.VT2 avdd 5.50471f
C123 a_28607_n287397# x2.delayPulse_digital_0/sky130_fd_sc_ls__xor2_1_0.X 0.190301f
C124 avdd x2.porPre 0.386243f
C125 a_30447_n288420# a_31045_n288085# 0.066235f
C126 avss a_17790_n286374# 0.045688f
C127 a_20598_n286374# a_21066_n286374# 0.307869f
C128 x2.delayPulse_digital_0/sky130_fd_sc_ls__xor2_1_0.X a_29214_n287320# 0.016368f
C129 a_14638_n288829# a_14970_n288829# 0.305459f
C130 w_31992_n290497# dvdd 1.0538f
C131 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N a_28056_n288420# 0.882223f
C132 x1.VD x1.Vinn 2.6259f
C133 x2.VT2 a_29876_n288037# 0.032579f
C134 a_21768_n288774# a_22236_n288774# 0.309677f
C135 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N a_28768_n287754# 0.012465f
C136 a_21534_n286374# avdd 0.112047f
C137 a_29688_n287709# a_29895_n287373# 0.220056f
C138 x1.vbn x1.VY 0.828345f
C139 a_21768_n288774# dvdd 0.041197f
C140 a_18259_n292308# a_18727_n292308# 0.309071f
C141 a_30447_n287429# dvdd 0.372127f
C142 a_13030_n290763# x1.vt 0.514642f
C143 a_19195_n292308# a_18727_n292308# 0.309071f
C144 a_29481_n287384# dvdd 0.385996f
C145 a_9762_n292173# x1.VD 0.768527f
C146 x1.VS a_13030_n290763# 0.758867f
C147 avss a_7606_n288829# 0.601486f
C148 a_19195_n292308# a_19663_n292308# 0.309071f
C149 a_10594_n288829# x1.Vinn 0.116674f
C150 a_10926_n288829# a_11258_n288829# 0.307869f
C151 avss a_13974_n288829# 0.334979f
C152 avdd x1.VY 0.795046f
C153 avss a_8822_n290308# 0.572442f
C154 x2.din avdd 1.17875f
C155 a_8436_n286429# a_8768_n286429# 0.307869f
C156 a_13642_n288829# x1.vt 0.118849f
C157 avss x1.vbn 10.528901f
C158 a_30814_n289746# x2.VT2 0.746546f
C159 x2.VT3 x1.vbn 0.016968f
C160 a_31045_n288085# x2.porPre 0.292728f
C161 avdd w_15901_n291463# 1.25112f
C162 avss avdd 43.161697f
C163 x2.VT3 avdd 1.71357f
C164 a_35074_n291454# x2.porPre 0.522625f
C165 x1.VY x1.Vinn 1.07195f
C166 a_18960_n288774# a_19428_n288774# 0.309677f
C167 a_35089_n289052# dvdd 1.56392f
C168 a_22002_n286374# a_22470_n286374# 0.307869f
C169 avss a_10428_n286429# 0.197326f
C170 a_32248_n290278# w_31992_n290497# 1.08624f
C171 x2.din a_15914_n289870# 1.20061f
C172 x2.x3.S1 avdd 0.114534f
C173 x2.Td_L a_28056_n288420# 0.05245f
C174 avdd a_30779_n287655# 0.032689f
C175 a_18493_n289908# a_18961_n289908# 0.309071f
C176 x1.VS x1.vt 0.180954f
C177 x1.VY a_9762_n292173# 1.1911f
C178 a_30022_n287538# dvdd 0.239037f
C179 a_19429_n289908# a_18961_n289908# 0.309071f
C180 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtp_1_0.D a_28607_n287397# 0.034956f
C181 x1.VD x1.Vinp 0.346443f
C182 a_19429_n289908# a_19897_n289908# 0.309071f
C183 a_11092_n286429# a_11424_n286429# 0.307869f
C184 x2.Td_L a_28768_n287754# 0.014868f
C185 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtp_1_0.D a_29214_n287320# 0.182152f
C186 w_15901_n291463# a_15914_n289870# 0.146582f
C187 a_19896_n288774# x2.din 0.045459f
C188 avss x1.Vinn 5.63805f
C189 a_20598_n286374# avdd 0.110373f
C190 x2.din a_20365_n289908# 0.042963f
C191 avss a_15914_n289870# 1.43798f
C192 a_20832_n288774# dvdd 0.041197f
C193 a_18727_n292308# vbg 0.05381f
C194 a_19663_n292308# vbg 0.05381f
C195 avss a_9100_n286429# 0.197326f
C196 a_23173_n289908# avdd 0.217187f
C197 x2.vbp1 dvdd 65.3681f
C198 avss a_9762_n292173# 0.606733f
C199 avdd x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A 8.12949f
C200 avss a_13144_n286429# 0.202195f
C201 a_30814_n289746# x2.VT3 0.170271f
C202 x1.vbn a_13030_n290763# 0.01692f
C203 a_19194_n286374# a_19662_n286374# 0.307869f
C204 a_21300_n288774# x2.din 0.045459f
C205 a_13642_n288829# a_13974_n288829# 0.309907f
C206 a_21067_n292308# a_21535_n292308# 0.309071f
C207 a_30410_n291353# w_31992_n290497# 0.063577f
C208 a_22002_n286374# avdd 0.117169f
C209 a_22236_n288774# dvdd 0.041197f
C210 avdd a_31115_n287366# 0.02289f
C211 avdd a_29688_n287709# 0.043511f
C212 avdd a_13030_n290763# 0.971935f
C213 a_28571_n287754# dvdd 0.010063f
C214 x2.x3.S1B dvdd 0.676749f
C215 a_8490_n290308# a_8822_n290308# 0.320088f
C216 avss a_7938_n288829# 0.335767f
C217 x1.VY x1.Vinp 0.383841f
C218 x2.VT2 porb_h[1] 0.317284f
C219 a_10926_n288829# x1.Vinn 0.116674f
C220 a_29487_n288398# dvdd 0.770655f
C221 a_29211_n288416# a_29671_n288104# 0.268084f
C222 avss a_14306_n288829# 0.334603f
C223 x2.porbPre x2.porPre 1.41505f
C224 x2.Td_S dvdd 2.17487f
C225 x2.vbp1 a_30112_n289746# 0.569749f
C226 x2.Td_L avdd 1.30208f
C227 a_7996_n292010# x1.VY 0.014688f
C228 avss a_17791_n292308# 0.046299f
C229 a_9930_n288829# a_10262_n288829# 0.307869f
C230 a_13974_n288829# x1.vt 0.118424f
C231 a_17790_n288774# dvdd 0.041943f
C232 avss x1.Vinp 6.34664f
C233 a_12978_n288829# a_12646_n288829# 0.312665f
C234 x2.VT2 porb_h[0] 0.15078f
C235 x2.VT2 w_31992_n290497# 0.324683f
C236 x2.delayPulse_digital_0/sky130_fd_sc_ls__xor2_1_0.X dvdd 0.583693f
C237 avss a_7996_n292010# 1.40406f
C238 x1.vbn x1.vt 0.052035f
C239 x1.vbn x1.VS 0.680843f
C240 a_30112_n289746# dvdd 1.06227f
C241 x2.Td_Lb dvdd 2.17504f
C242 x2.Td_Lb a_29487_n288398# 0.251149f
C243 a_13808_n286429# a_14140_n286429# 0.309907f
C244 a_21301_n289908# a_21769_n289908# 0.309071f
C245 avss a_10760_n286429# 0.197326f
C246 avdd a_29895_n287373# 0.026079f
C247 x2.VT2 a_30447_n287429# 0.014496f
C248 x2.VT2 a_29481_n287384# 0.017194f
C249 avdd x1.vt 7.16197f
C250 avdd x1.VS 1.0014f
C251 avdd a_29211_n288416# 0.014059f
C252 a_30011_n288135# dvdd 0.202587f
C253 a_29487_n288398# a_30011_n288135# 0.049973f
C254 a_20364_n288774# x2.din 0.045459f
C255 a_21066_n286374# avdd 0.111083f
C256 x2.din a_20833_n289908# 0.042963f
C257 a_10096_n286429# a_10428_n286429# 0.307869f
C258 a_28607_n287397# x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N 0.021397f
C259 a_32248_n290278# dvdd 1.25433f
C260 a_20131_n292308# vbg 0.05381f
C261 avss a_9432_n286429# 0.197326f
C262 a_29211_n288416# a_29876_n288037# 0.195254f
C263 a_8602_n288829# a_8934_n288829# 0.307869f
C264 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N a_29214_n287320# 0.039522f
C265 a_18024_n288774# dvdd 0.045757f
C266 x1.vt x1.Vinn 0.023838f
C267 x2.porbPre x2.x3.S1 0.547836f
C268 a_13144_n286429# a_12812_n286429# 0.312665f
C269 x2.vbp1 por 0.581019f
C270 x1.VS x1.Vinn 1.09827f
C271 x1.vt a_15914_n289870# 0.212492f
C272 x2.vbp1 x2.x3.aout 0.031103f
C273 avss a_13476_n286429# 0.201521f
C274 a_21768_n288774# x2.din 0.045459f
C275 a_22236_n288774# a_22704_n288774# 0.309677f
C276 avdd a_17790_n286374# 0.112582f
C277 x2.Td_Lb a_30011_n288135# 0.152772f
C278 x1.VS a_9762_n292173# 0.416229f
C279 a_13030_n290763# x1.Vinp 0.697845f
C280 x2.VT3 w_31992_n290497# 1.75603f
C281 a_22470_n286374# avdd 0.414269f
C282 a_22704_n288774# dvdd 0.041197f
C283 a_17790_n288774# a_18024_n288774# 0.311625f
C284 x2.VT2 a_30022_n287538# 0.043926f
C285 avss a_8270_n288829# 0.335767f
C286 avdd a_29671_n288104# 0.03834f
C287 a_19663_n292308# a_20131_n292308# 0.309071f
C288 a_30447_n288420# dvdd 0.368159f
C289 a_29487_n288398# a_30447_n288420# 0.034318f
C290 a_11258_n288829# x1.Vinn 0.424902f
C291 a_29671_n288104# a_30699_n288291# 0.078258f
C292 avss a_14638_n288829# 0.335276f
C293 dvdd por 8.63071f
C294 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A porb_h[1] 3.00808f
C295 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtp_1_0.D dvdd 1.42566f
C296 a_18258_n286374# a_17790_n286374# 0.307869f
C297 x2.x3.aout dvdd 0.310939f
C298 x1.Vinp a_12812_n286429# 0.316525f
C299 a_29671_n288104# a_29876_n288037# 0.098669f
C300 a_14306_n288829# x1.vt 0.117999f
C301 a_8768_n286429# a_9100_n286429# 0.307869f
C302 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N a_29481_n287384# 0.174319f
C303 x2.vbp1 x2.VT2 0.068045f
C304 a_30779_n287655# a_30447_n287429# 0.251184f
C305 a_29481_n287384# a_30779_n287655# 0.058581f
C306 a_29214_n287320# a_29688_n287709# 0.314195f
C307 x2.porbPre a_31115_n287366# 0.087517f
C308 x2.Td_L a_28607_n287397# 0.096203f
C309 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A porb_h[0] 2.88344f
C310 x2.vbp2 avdd 0.432735f
C311 avdd x1.vbn 0.72255f
C312 a_19428_n288774# a_19896_n288774# 0.309677f
C313 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtp_1_0.D x2.delayPulse_digital_0/sky130_fd_sc_ls__xor2_1_0.X 0.385496f
C314 a_22470_n286374# a_22938_n286374# 0.307869f
C315 x2.Td_Lb a_30447_n288420# 0.262864f
C316 avss a_12646_n288829# 0.499575f
C317 x1.vt x1.Vinp 0.044922f
C318 x1.VS x1.Vinp 1.22558f
C319 avss a_11092_n286429# 0.197326f
C320 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtp_1_0.D x2.Td_Lb 0.228134f
C321 avdd a_30699_n288291# 0.036749f
C322 a_19897_n289908# a_20365_n289908# 0.309071f
C323 x2.VT2 dvdd 2.67927f
C324 x2.porPre dvdd 1.7449f
C325 a_30011_n288135# a_30447_n288420# 0.16939f
C326 a_20832_n288774# x2.din 0.045459f
C327 x2.din a_21301_n289908# 0.042963f
C328 x2.Td_L w_31992_n290497# 0.057323f
C329 avdd a_29876_n288037# 0.03731f
C330 a_20599_n292308# vbg 0.05381f
C331 avss a_9764_n286429# 0.197326f
C332 avss a_9930_n288829# 0.329279f
C333 a_18258_n286374# avdd 0.110373f
C334 a_30447_n287429# a_31115_n287366# 0.083162f
C335 a_29688_n287709# a_30447_n287429# 0.153568f
C336 a_29214_n287320# a_29895_n287373# 0.045318f
C337 a_29481_n287384# a_29688_n287709# 0.418019f
C338 a_18492_n288774# dvdd 0.042912f
C339 x1.vbn a_9762_n292173# 0.084991f
C340 avdd x1.Vinn 0.710534f
C341 avdd a_15914_n289870# 0.339476f
C342 avss vbg 11.2283f
C343 a_7606_n288829# a_7938_n288829# 0.307869f
C344 x2.VT3 vbg 0.026316f
C345 avss a_13808_n286429# 0.200846f
C346 x2.vbp2 a_30814_n289746# 0.338088f
C347 a_30112_n289746# x2.VT2 0.081907f
C348 x2.vbp1 x2.VT3 1.40074f
C349 a_19662_n286374# a_20130_n286374# 0.307869f
C350 x2.VT2 x2.Td_Lb 0.131131f
C351 a_22236_n288774# x2.din 0.045459f
C352 x2.Td_Lb x2.porPre 0.801193f
C353 a_21535_n292308# a_22003_n292308# 0.309071f
C354 a_13974_n288829# a_14306_n288829# 0.309029f
C355 avdd a_9762_n292173# 0.677366f
C356 a_22938_n286374# avdd 0.630465f
C357 x2.din dvdd 2.31677f
C358 a_30814_n289746# avdd 0.584939f
C359 avss a_8602_n288829# 0.335767f
C360 avdd a_31045_n288085# 0.029777f
C361 x2.VT2 a_30011_n288135# 0.030428f
C362 a_30699_n288291# a_31045_n288085# 0.076493f
C363 avss a_14970_n288829# 1.5487f
C364 a_17790_n288774# a_18025_n289908# 0.309983f
C365 a_10262_n288829# a_10594_n288829# 0.307869f
C366 x2.VT2 a_32248_n290278# 0.039716f
C367 avss dvdd 1.28718f
C368 a_23173_n289908# vbg 0.573644f
C369 x2.VT3 dvdd 0.7414f
C370 a_17790_n288774# x2.din 0.369627f
C371 a_14638_n288829# x1.vt 0.118923f
C372 a_28607_n287397# a_28768_n287754# 0.190208f
C373 x2.x3.S1 x2.x3.S1B 1.1152f
C374 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N dvdd 1.09002f
C375 x2.x3.S1 dvdd 1.56456f
C376 a_29481_n287384# a_29895_n287373# 0.070205f
C377 a_29688_n287709# a_30022_n287538# 0.314482f
C378 x2.vbp1 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A 0.054194f
C379 a_30779_n287655# dvdd 0.305597f
C380 a_7772_n286429# a_8104_n286429# 0.307869f
C381 x1.vbn a_7996_n292010# 0.685806f
C382 a_17790_n288774# avss 0.063911f
C383 a_21769_n289908# a_22237_n289908# 0.309071f
C384 a_14140_n286429# a_14472_n286429# 0.309029f
C385 avss a_8656_n292108# 0.596837f
C386 avdd x1.Vinp 0.442449f
C387 avss a_11424_n286429# 0.381741f
C388 a_9930_n288829# a_9598_n288829# 0.307869f
C389 a_18024_n288774# a_18492_n288774# 0.309677f
C390 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N x2.delayPulse_digital_0/sky130_fd_sc_ls__xor2_1_0.X 0.095428f
C391 x2.VT2 a_30447_n288420# 0.017933f
C392 x2.VT3 x2.Td_Lb 0.017295f
C393 a_18024_n288774# a_18025_n289908# 0.021824f
C394 a_30447_n288420# x2.porPre 0.011381f
C395 avdd porb 0.199778f
C396 x1.vt a_12646_n288829# 0.017673f
C397 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A dvdd 0.6058f
C398 x2.din a_21769_n289908# 0.042963f
C399 x2.VT2 a_30410_n291353# 0.580175f
C400 a_10428_n286429# a_10760_n286429# 0.307869f
C401 a_21067_n292308# vbg 0.05381f
C402 a_18024_n288774# x2.din 0.012958f
C403 x1.Vinn x1.Vinp 1.95521f
C404 a_8934_n288829# a_9266_n288829# 0.307869f
C405 a_27214_n288191# dvdd 1.11143f
C406 a_22471_n292308# a_22003_n292308# 0.309071f
C407 avss a_10262_n288829# 0.306053f
C408 a_18726_n286374# avdd 0.110373f
C409 a_30022_n287538# a_29895_n287373# 0.260781f
C410 a_18960_n288774# dvdd 0.041422f
C411 a_31115_n287366# dvdd 0.261137f
C412 a_29688_n287709# dvdd 0.168597f
C413 x2.VT3 a_32248_n290278# 0.388549f
C414 avss a_7772_n286429# 0.505195f
C415 avdd porb_h[1] 4.47236f
C416 x2.porbPre avdd 0.384944f
C417 avss a_14140_n286429# 0.20017f
C418 a_22704_n288774# x2.din 0.045569f
C419 x2.Td_L dvdd 4.24551f
C420 a_10096_n286429# a_9764_n286429# 0.307869f
C421 x2.vbp2 w_31992_n290497# 0.398779f
C422 a_18258_n286374# a_18726_n286374# 0.307869f
C423 avss a_8934_n288829# 0.335767f
C424 a_12978_n288829# a_13310_n288829# 0.311725f
C425 a_20131_n292308# a_20599_n292308# 0.309071f
C426 avdd porb_h[0] 4.4046f
C427 avdd w_31992_n290497# 1.67875f
C428 avss a_12978_n288829# 0.337152f
C429 x2.Td_L x2.delayPulse_digital_0/sky130_fd_sc_ls__xor2_1_0.X 0.296806f
C430 a_14970_n288829# x1.vt 0.315571f
C431 a_9100_n286429# a_9432_n286429# 0.307869f
C432 a_22705_n289908# a_22237_n289908# 0.309071f
C433 x2.Td_L x2.Td_Lb 3.39981f
C434 avdd a_30447_n287429# 0.059189f
C435 avdd a_29481_n287384# 0.033726f
C436 x1.VY x1.VD 2.11152f
C437 a_29895_n287373# dvdd 0.325593f
C438 a_29895_n287373# a_29487_n288398# 0.01331f
C439 x2.VT3 a_30410_n291353# 0.894634f
C440 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtp_1_0.D x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N 0.388955f
C441 x1.vt dvdd 0.036968f
C442 a_29211_n288416# dvdd 0.313389f
C443 a_29211_n288416# a_29487_n288398# 0.123863f
C444 a_19896_n288774# a_20364_n288774# 0.309677f
C445 x2.din a_22705_n289908# 0.042963f
C446 a_13144_n286429# a_13476_n286429# 0.311725f
C447 a_20365_n289908# a_20833_n289908# 0.309071f
C448 a_22471_n292308# a_22939_n292308# 0.309071f
C449 avss x1.VD 3.02338f
C450 a_30814_n289746# w_31992_n290497# 0.096314f
C451 x2.din a_22237_n289908# 0.042963f
C452 x2.VT2 avss 0.138801f
C453 x2.VT2 x2.VT3 1.17092f
C454 a_21535_n292308# vbg 0.05381f
C455 a_18492_n288774# x2.din 0.052229f
C456 a_28056_n288420# dvdd 0.874706f
C457 x2.Td_Lb a_29211_n288416# 0.251053f
C458 avss a_10594_n288829# 0.239853f
C459 x2.din a_18025_n289908# 0.012607f
C460 a_19194_n286374# avdd 0.110373f
C461 a_19428_n288774# dvdd 0.041197f
C462 a_27214_n288191# x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtp_1_0.D 0.239718f
C463 avdd a_30022_n287538# 0.042554f
C464 a_28768_n287754# dvdd 0.19655f
C465 avss a_8104_n286429# 0.197326f
C466 a_7938_n288829# a_8270_n288829# 0.307869f
C467 x1.vbn vbg 0.015171f
C468 a_29671_n288104# dvdd 0.22226f
C469 a_29487_n288398# a_29671_n288104# 0.469956f
C470 avss a_14472_n286429# 0.199494f
C471 a_20130_n286374# a_20598_n286374# 0.307869f
C472 x2.vbp1 x2.vbp2 0.809231f
C473 a_14306_n288829# a_14638_n288829# 0.308171f
C474 a_20598_n286374# x2.VT2 0.011586f
C475 x2.delayPulse_digital_0/sky130_fd_sc_ls__xor2_1_0.X a_28056_n288420# 0.487997f
C476 avdd vbg 8.42169f
C477 x2.Td_L x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtp_1_0.D 0.043867f
C478 a_21300_n288774# a_21768_n288774# 0.309677f
C479 avss a_9266_n288829# 0.335767f
C480 x2.vbp1 avdd 0.966462f
C481 a_22705_n289908# a_23173_n289908# 0.309071f
C482 avss x1.VY 2.28271f
C483 x2.delayPulse_digital_0/sky130_fd_sc_ls__xor2_1_0.X a_28768_n287754# 0.062836f
C484 x2.VT2 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A 0.452889f
C485 a_17791_n292308# a_18259_n292308# 0.309071f
C486 x2.din avss 1.24529f
C487 a_10594_n288829# a_10926_n288829# 0.307869f
C488 avss a_13310_n288829# 0.336926f
C489 x2.VT3 a_20599_n292308# 0.010992f
C490 por dvss 5.558747f
C491 vbg dvss 26.75568f
C492 porb dvss 6.743152f
C493 porb_h[1] dvss 3.891496f
C494 porb_h[0] dvss 4.959771f
C495 dvdd dvss 0.101262p
C496 avdd dvss 0.296748p
C497 avss dvss 67.802795f
C498 a_35074_n291454# dvss 0.98581f
C499 a_30410_n291353# dvss 2.10904f
C500 a_32248_n290278# dvss 1.592f
C501 a_25216_n290828# dvss 0.250795f
C502 x2.VT3 dvss 1.01851p
C503 x2.VT2 dvss 1.024111p
C504 a_30814_n289746# dvss 0.050779f
C505 x2.vbp2 dvss 1.14188f
C506 a_30112_n289746# dvss 0.079624f
C507 x2.vbp1 dvss 18.344463f
C508 a_23173_n289908# dvss 7.24083f
C509 a_22939_n292308# dvss 1.05749f
C510 a_22705_n289908# dvss 0.736313f
C511 a_22471_n292308# dvss 0.744182f
C512 a_22237_n289908# dvss 0.659075f
C513 a_22003_n292308# dvss 0.724196f
C514 a_21769_n289908# dvss 0.77106f
C515 a_21535_n292308# dvss 0.712586f
C516 a_21301_n289908# dvss 0.771552f
C517 a_21067_n292308# dvss 0.707345f
C518 a_20833_n289908# dvss 0.771552f
C519 a_20599_n292308# dvss 0.712197f
C520 a_20365_n289908# dvss 0.771552f
C521 a_20131_n292308# dvss 0.712302f
C522 a_19897_n289908# dvss 0.771552f
C523 a_19663_n292308# dvss 0.712302f
C524 a_19429_n289908# dvss 0.771552f
C525 a_19195_n292308# dvss 0.712561f
C526 a_18961_n289908# dvss 0.759035f
C527 a_18727_n292308# dvss 0.714044f
C528 a_18493_n289908# dvss 0.742346f
C529 a_18259_n292308# dvss 0.714974f
C530 a_18025_n289908# dvss 0.723692f
C531 a_17791_n292308# dvss 0.948058f
C532 a_15914_n289870# dvss 0.501302f
C533 x1.vt dvss 1.918339f
C534 a_13030_n290763# dvss 0.274602f
C535 x1.VD dvss 4.241671f
C536 a_9762_n292173# dvss 0.327888f
C537 x1.VS dvss 1.71665f
C538 x1.VY dvss 3.296263f
C539 a_8822_n290308# dvss 0.153358f
C540 a_8656_n292108# dvss 0.2732f
C541 a_8490_n290308# dvss 0.154081f
C542 a_7996_n292010# dvss 0.658692f
C543 x1.vbn dvss 7.085366f
C544 a_35089_n289052# dvss 0.889652f
C545 a_29876_n288037# dvss 0.21181f
C546 x2.porPre dvss 2.93939f
C547 a_31045_n288085# dvss 0.358048f
C548 a_30447_n288420# dvss 0.41534f
C549 a_30699_n288291# dvss 0.37154f
C550 a_30011_n288135# dvss 0.18597f
C551 a_29671_n288104# dvss 1.11242f
C552 a_29487_n288398# dvss 0.629109f
C553 a_29211_n288416# dvss 0.225211f
C554 x2.Td_Lb dvss 4.36387f
C555 a_28056_n288420# dvss 1.41269f
C556 a_28768_n287754# dvss 0.012546f
C557 a_31115_n287366# dvss 0.295369f
C558 a_30447_n287429# dvss 0.576108f
C559 a_30779_n287655# dvss 0.213838f
C560 x2.x3.aout dvss 2.567305f
C561 x2.x3.S1B dvss 2.34613f
C562 a_29895_n287373# dvss 0.134629f
C563 a_30022_n287538# dvss 0.172993f
C564 a_29688_n287709# dvss 0.985543f
C565 a_29481_n287384# dvss 1.12579f
C566 a_29214_n287320# dvss 0.31512f
C567 x2.delayPulse_digital_0/sky130_fd_sc_ls__xor2_1_0.X dvss 1.90063f
C568 a_28868_n287397# dvss 0.01266f
C569 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.CLK_N dvss 1.49183f
C570 a_28607_n287397# dvss 0.301715f
C571 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtp_1_0.D dvss 2.23981f
C572 a_27214_n288191# dvss 1.72706f
C573 x2.Td_L dvss 5.218703f
C574 x2.x3.S1 dvss 3.31642f
C575 x2.porbPre dvss 3.80558f
C576 x2.Td_S dvss 2.58821f
C577 x2.din dvss 8.02483f
C578 a_22938_n286374# dvss 0.857375f
C579 a_22704_n288774# dvss 0.909569f
C580 a_22470_n286374# dvss 0.657786f
C581 a_22236_n288774# dvss 0.641564f
C582 a_22002_n286374# dvss 0.702374f
C583 a_21768_n288774# dvss 0.769918f
C584 a_21534_n286374# dvss 0.703445f
C585 a_21300_n288774# dvss 0.770175f
C586 a_21066_n286374# dvss 0.702533f
C587 a_20832_n288774# dvss 0.770174f
C588 a_20598_n286374# dvss 0.706444f
C589 a_20364_n288774# dvss 0.770174f
C590 a_20130_n286374# dvss 0.703445f
C591 a_19896_n288774# dvss 0.770174f
C592 a_19662_n286374# dvss 0.703445f
C593 a_19428_n288774# dvss 0.770272f
C594 a_19194_n286374# dvss 0.703445f
C595 a_18960_n288774# dvss 0.755679f
C596 a_18726_n286374# dvss 0.703445f
C597 a_18492_n288774# dvss 0.741396f
C598 a_18258_n286374# dvss 0.700806f
C599 a_18024_n288774# dvss 0.720897f
C600 a_17790_n288774# dvss 1.52514f
C601 a_17790_n286374# dvss 0.893304f
C602 a_14970_n288829# dvss 0.175412f
C603 a_14804_n286429# dvss 0.362007f
C604 a_14638_n288829# dvss 0.241028f
C605 a_14472_n286429# dvss 0.361214f
C606 a_14306_n288829# dvss 0.241024f
C607 a_14140_n286429# dvss 0.361588f
C608 a_13974_n288829# dvss 0.240951f
C609 a_13808_n286429# dvss 0.36743f
C610 a_13642_n288829# dvss 0.240877f
C611 a_13476_n286429# dvss 0.356698f
C612 a_13310_n288829# dvss 0.240803f
C613 a_13144_n286429# dvss 0.36271f
C614 a_12978_n288829# dvss 0.24073f
C615 a_12812_n286429# dvss 0.362653f
C616 a_12646_n288829# dvss 0.240652f
C617 x1.Vinp dvss 2.733891f
C618 x1.Vinn dvss 2.246496f
C619 a_11424_n286429# dvss 0.388305f
C620 a_11258_n288829# dvss 0.240962f
C621 a_11092_n286429# dvss 0.36015f
C622 a_10926_n288829# dvss 0.240962f
C623 a_10760_n286429# dvss 0.36015f
C624 a_10594_n288829# dvss 0.240962f
C625 a_10428_n286429# dvss 0.356539f
C626 a_10262_n288829# dvss 0.240962f
C627 a_10096_n286429# dvss 0.37682f
C628 a_9930_n288829# dvss 0.240962f
C629 a_9764_n286429# dvss 0.354717f
C630 a_9598_n288829# dvss 0.240962f
C631 a_9432_n286429# dvss 0.36015f
C632 a_9266_n288829# dvss 0.240962f
C633 a_9100_n286429# dvss 0.36015f
C634 a_8934_n288829# dvss 0.240962f
C635 a_8768_n286429# dvss 0.36015f
C636 a_8602_n288829# dvss 0.240962f
C637 a_8436_n286429# dvss 0.36015f
C638 a_8270_n288829# dvss 0.240962f
C639 a_8104_n286429# dvss 0.36015f
C640 a_7938_n288829# dvss 0.240962f
C641 a_7772_n286429# dvss 0.36015f
C642 a_7606_n288829# dvss 0.240962f
C643 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A dvss 13.209143f
C644 w_31992_n290497# dvss 2.3241f
C645 w_15901_n291463# dvss 1.98573f
C646 vbg.t0 dvss 0.81819f
C647 x1.VY.n0 dvss 0.489423f
C648 x1.VY.t0 dvss 0.080438f
C649 x1.VY.t2 dvss 0.038968f
C650 x1.VY.t3 dvss 0.081006f
C651 x1.VY.t1 dvss 0.03921f
C652 x1.VY.t5 dvss 0.112609f
C653 x1.VY.t4 dvss 0.086221f
C654 x1.VY.t6 dvss 0.082418f
C655 x1.VY.n1 dvss 1.28976f
C656 x1.vo1.n0 dvss 1.23665f
C657 x1.x1.S dvss 1.5909f
C658 x1.vo1.t8 dvss 0.214756f
C659 x1.vo1.t4 dvss 0.213887f
C660 x1.vo1.n1 dvss 0.592208f
C661 x1.vo1.t1 dvss 0.071042f
C662 x1.vo1.t5 dvss 0.212934f
C663 x1.vo1.t3 dvss 0.207223f
C664 x1.vo1.t7 dvss 0.30217f
C665 x1.vo1.t6 dvss 0.317878f
C666 x1.vo1.t2 dvss 0.214917f
C667 x1.vo1.n2 dvss 0.980634f
C668 x1.vo1.t0 dvss 0.271722f
C669 x1.vo1.n3 dvss 1.77308f
C670 a_4566_n290308.t1 dvss 2.20295f
C671 a_4566_n290308.t0 dvss 0.048713f
C672 a_4566_n290308.t2 dvss 0.048336f
C673 a_4508_n291419.t0 dvss 1.9171f
C674 a_4508_n291419.t2 dvss 0.041648f
C675 a_4508_n291419.t1 dvss 0.041254f
C676 x1.Vinp.t3 dvss 0.539496f
C677 x1.Vinp.t2 dvss 0.538514f
C678 x1.Vinp.n0 dvss 1.2311f
C679 x1.Vinp.t0 dvss 0.064016f
C680 x1.Vinp.t1 dvss 0.064175f
C681 x1.Vinp.n1 dvss 2.31708f
C682 a_24570_n290925.n0 dvss 0.516596f
C683 a_24570_n290925.t0 dvss 13.4951f
C684 a_24570_n290925.t2 dvss 0.124375f
C685 a_24570_n290925.t4 dvss 0.12543f
C686 a_24570_n290925.t1 dvss 0.021863f
C687 a_24570_n290925.n1 dvss 1.47877f
C688 a_24570_n290925.t3 dvss 0.037901f
C689 x2.Td_S.n0 dvss 0.782416f
C690 x2.Td_S.t0 dvss 0.036142f
C691 x2.Td_S.t5 dvss 0.059231f
C692 x2.Td_S.t6 dvss 0.061137f
C693 x2.Td_S.t4 dvss 0.059626f
C694 x2.Td_S.t3 dvss 0.072423f
C695 x2.Td_S.t2 dvss 0.071471f
C696 x2.Td_S.t1 dvss 0.036622f
C697 a_24253_n287224.n0 dvss 0.540224f
C698 a_24253_n287224.n1 dvss 2.7426f
C699 a_24253_n287224.n2 dvss 0.754469f
C700 a_24253_n287224.n3 dvss 0.372496f
C701 a_24253_n287224.t4 dvss 0.116416f
C702 a_24253_n287224.t11 dvss 0.116237f
C703 a_24253_n287224.t7 dvss 0.140184f
C704 a_24253_n287224.t5 dvss 0.139789f
C705 a_24253_n287224.n4 dvss 0.634023f
C706 a_24253_n287224.n5 dvss 1.88264f
C707 a_24253_n287224.t1 dvss 0.042178f
C708 a_24253_n287224.t0 dvss 0.042702f
C709 a_24253_n287224.t9 dvss 0.116149f
C710 a_24253_n287224.t6 dvss 0.115962f
C711 a_24253_n287224.t8 dvss 0.140375f
C712 a_24253_n287224.t10 dvss 0.13931f
C713 a_24253_n287224.t2 dvss 0.082121f
C714 a_24253_n287224.t3 dvss 0.082121f
C715 x1.VD.n0 dvss 1.9551f
C716 x1.VD.n1 dvss 1.84602f
C717 x1.VD.t2 dvss 0.069792f
C718 x1.VD.t0 dvss 0.132548f
C719 x1.VD.n2 dvss 0.686392f
C720 x1.VD.t7 dvss 0.138045f
C721 x1.VD.t4 dvss 0.136638f
C722 x1.VD.t5 dvss 0.136333f
C723 x1.VD.t1 dvss 0.288665f
C724 x1.VD.n3 dvss 0.982727f
C725 x1.VD.t3 dvss 0.137072f
C726 x1.VD.t6 dvss 0.136839f
C727 x1.VD.t8 dvss 0.138216f
C728 x1.VD.n4 dvss 0.985802f
C729 x2.x3.aout.n0 dvss 1.38768f
C730 x2.x3.aout.n1 dvss 0.788589f
C731 x2.x3.aout.t3 dvss 0.17003f
C732 x2.x3.aout.t5 dvss 0.102937f
C733 x2.x3.aout.t4 dvss 0.17003f
C734 x2.x3.aout.t6 dvss 0.102937f
C735 x2.x3.aout.t0 dvss 0.064956f
C736 x2.x3.aout.t1 dvss 0.106636f
C737 x2.x3.aout.t2 dvss 0.106046f
C738 a_13449_n292106.t3 dvss 0.371455f
C739 a_13449_n292106.t1 dvss 0.3701f
C740 a_13449_n292106.t0 dvss 0.311387f
C741 a_13449_n292106.n0 dvss 2.1121f
C742 a_13449_n292106.t2 dvss 0.234955f
C743 x2.vbn1.n0 dvss 0.065145f
C744 x2.vbn1.n1 dvss 0.05439f
C745 x2.vbn1.t0 dvss 5.38468f
C746 x2.vbn1.t19 dvss 0.014905f
C747 x2.vbn1.t16 dvss 0.015058f
C748 x2.vbn1.n2 dvss 0.031655f
C749 x2.vbn1.t20 dvss 0.014905f
C750 x2.vbn1.t17 dvss 0.014905f
C751 x2.vbn1.t18 dvss 0.014905f
C752 x2.vbn1.t7 dvss 0.014905f
C753 x2.vbn1.t1 dvss 0.014905f
C754 x2.vbn1.t9 dvss 0.014905f
C755 x2.vbn1.t11 dvss 0.014905f
C756 x2.vbn1.t5 dvss 0.014905f
C757 x2.vbn1.t3 dvss 0.014905f
C758 x2.vbn1.t13 dvss 0.014905f
C759 x2.vbn1.n6 dvss 0.188857f
C760 x2.vbn1.n7 dvss 0.018158f
C761 x2.vbn1.n8 dvss 0.016268f
C762 x2.vbn1.n9 dvss 0.016272f
C763 x2.vbn1.n10 dvss 0.016264f
C764 x2.vbn1.n11 dvss 0.016264f
C765 x2.vbn1.n12 dvss 0.01629f
C766 x2.vbn1.n13 dvss 0.017297f
C767 x2.vbn1.n14 dvss 0.018333f
C768 x2.vbn1.n15 dvss 0.017345f
C769 x2.vbn1.n16 dvss 0.016272f
C770 a_34015_n286994.n0 dvss 1.10914f
C771 a_34015_n286994.n1 dvss 0.320385f
C772 a_34015_n286994.n2 dvss 0.195689f
C773 a_34015_n286994.t4 dvss 0.186945f
C774 a_34015_n286994.t5 dvss 0.186787f
C775 a_34015_n286994.n3 dvss 0.157412f
C776 a_34015_n286994.t2 dvss 0.108582f
C777 a_34015_n286994.t0 dvss 0.065409f
C778 a_34015_n286994.t1 dvss 0.065552f
C779 a_34015_n286994.t3 dvss 0.104095f
C780 a_24270_n290121.n0 dvss 2.20563f
C781 a_24270_n290121.n1 dvss 0.441814f
C782 a_24270_n290121.t0 dvss 49.9608f
C783 a_24270_n290121.t3 dvss 0.011213f
C784 a_24270_n290121.t5 dvss 0.011213f
C785 a_24270_n290121.t15 dvss 0.011213f
C786 a_24270_n290121.n2 dvss 0.024915f
C787 a_24270_n290121.t9 dvss 0.011213f
C788 a_24270_n290121.t17 dvss 0.011213f
C789 a_24270_n290121.n3 dvss 0.024198f
C790 a_24270_n290121.n4 dvss 0.419817f
C791 a_24270_n290121.t1 dvss 0.042317f
C792 a_24270_n290121.t6 dvss 0.134597f
C793 a_24270_n290121.t10 dvss 0.134597f
C794 a_24270_n290121.t12 dvss 0.134597f
C795 a_24270_n290121.t2 dvss 0.134597f
C796 a_24270_n290121.t16 dvss 0.134597f
C797 a_24270_n290121.t8 dvss 0.134597f
C798 a_24270_n290121.t18 dvss 0.135131f
C799 a_24270_n290121.t14 dvss 0.134597f
C800 a_24270_n290121.t4 dvss 0.135884f
C801 a_24270_n290121.n5 dvss 0.148815f
C802 a_24270_n290121.n6 dvss 0.15021f
C803 a_24270_n290121.n7 dvss 0.149959f
C804 a_24270_n290121.n8 dvss 0.149994f
C805 a_24270_n290121.n9 dvss 0.150102f
C806 a_24270_n290121.n10 dvss 0.166517f
C807 a_24270_n290121.t11 dvss 0.011213f
C808 a_24270_n290121.t7 dvss 0.011213f
C809 a_24270_n290121.n11 dvss 0.024188f
C810 a_24270_n290121.n12 dvss 0.219145f
C811 a_24270_n290121.n13 dvss 0.194509f
C812 a_24270_n290121.n14 dvss 0.024219f
C813 a_24270_n290121.t13 dvss 0.011213f
C814 x1.Vinn.t2 dvss 0.443587f
C815 x1.Vinn.t6 dvss 0.442708f
C816 x1.Vinn.n0 dvss 0.83768f
C817 x1.Vinn.t3 dvss 0.443578f
C818 x1.Vinn.t7 dvss 0.442706f
C819 x1.Vinn.n1 dvss 0.78681f
C820 x1.Vinn.n2 dvss 0.210885f
C821 x1.Vinn.t4 dvss 0.442715f
C822 x1.Vinn.t5 dvss 0.443655f
C823 x1.Vinn.n3 dvss 0.783772f
C824 x1.Vinn.n4 dvss 0.132744f
C825 x1.Vinn.t1 dvss 0.053095f
C826 x1.Vinn.t0 dvss 0.236839f
C827 x1.Vinn.n5 dvss 1.56633f
C828 a_35277_n289052.t2 dvss 0.014535f
C829 a_35277_n289052.t1 dvss 0.010382f
C830 a_35277_n289052.t0 dvss 0.010382f
C831 a_35277_n289052.n0 dvss 0.023071f
C832 a_35277_n289052.t9 dvss 0.011326f
C833 a_35277_n289052.t25 dvss 0.011326f
C834 a_35277_n289052.t29 dvss 0.011326f
C835 a_35277_n289052.t17 dvss 0.023763f
C836 a_35277_n289052.n1 dvss 0.067184f
C837 a_35277_n289052.n2 dvss 0.046663f
C838 a_35277_n289052.n3 dvss 0.036696f
C839 a_35277_n289052.t18 dvss 0.011326f
C840 a_35277_n289052.t27 dvss 0.011326f
C841 a_35277_n289052.t13 dvss 0.011326f
C842 a_35277_n289052.t23 dvss 0.023763f
C843 a_35277_n289052.n4 dvss 0.067184f
C844 a_35277_n289052.n5 dvss 0.046663f
C845 a_35277_n289052.n6 dvss 0.036696f
C846 a_35277_n289052.n7 dvss 0.055758f
C847 a_35277_n289052.t11 dvss 0.028126f
C848 a_35277_n289052.t21 dvss 0.030297f
C849 a_35277_n289052.t24 dvss 0.028126f
C850 a_35277_n289052.t12 dvss 0.030297f
C851 a_35277_n289052.t6 dvss 0.028126f
C852 a_35277_n289052.t16 dvss 0.030297f
C853 a_35277_n289052.t19 dvss 0.028126f
C854 a_35277_n289052.t7 dvss 0.041066f
C855 a_35277_n289052.n8 dvss 0.074326f
C856 a_35277_n289052.n9 dvss 0.0494f
C857 a_35277_n289052.n10 dvss 0.039433f
C858 a_35277_n289052.t20 dvss 0.028126f
C859 a_35277_n289052.t8 dvss 0.030297f
C860 a_35277_n289052.t28 dvss 0.028126f
C861 a_35277_n289052.t15 dvss 0.030297f
C862 a_35277_n289052.t14 dvss 0.028126f
C863 a_35277_n289052.t26 dvss 0.030297f
C864 a_35277_n289052.t22 dvss 0.028126f
C865 a_35277_n289052.t10 dvss 0.041066f
C866 a_35277_n289052.n11 dvss 0.074326f
C867 a_35277_n289052.n12 dvss 0.0494f
C868 a_35277_n289052.n13 dvss 0.039433f
C869 a_35277_n289052.n14 dvss 0.054971f
C870 a_35277_n289052.n15 dvss 0.77802f
C871 a_35277_n289052.n16 dvss 0.309365f
C872 a_35277_n289052.t4 dvss 0.014535f
C873 a_35277_n289052.t3 dvss 0.014535f
C874 a_35277_n289052.n17 dvss 0.030267f
C875 a_35277_n289052.n18 dvss 0.30772f
C876 a_35277_n289052.n19 dvss 0.030112f
C877 a_35277_n289052.t5 dvss 0.014535f
C878 porb.t7 dvss 0.018111f
C879 porb.t0 dvss 0.018111f
C880 porb.n0 dvss 0.040123f
C881 porb.t28 dvss 0.025356f
C882 porb.t16 dvss 0.025356f
C883 porb.n1 dvss 0.0528f
C884 porb.t45 dvss 0.025356f
C885 porb.t33 dvss 0.025356f
C886 porb.n2 dvss 0.052529f
C887 porb.n3 dvss 0.521914f
C888 porb.t10 dvss 0.018111f
C889 porb.t4 dvss 0.018111f
C890 porb.n4 dvss 0.040174f
C891 porb.t35 dvss 0.025356f
C892 porb.t25 dvss 0.025356f
C893 porb.n5 dvss 0.0528f
C894 porb.t21 dvss 0.025356f
C895 porb.t42 dvss 0.025356f
C896 porb.n6 dvss 0.052529f
C897 porb.n7 dvss 0.52367f
C898 porb.t14 dvss 0.018111f
C899 porb.t8 dvss 0.018111f
C900 porb.n8 dvss 0.040174f
C901 porb.t43 dvss 0.025356f
C902 porb.t30 dvss 0.025356f
C903 porb.n9 dvss 0.0528f
C904 porb.t29 dvss 0.025356f
C905 porb.t47 dvss 0.025356f
C906 porb.n10 dvss 0.052529f
C907 porb.n11 dvss 0.52367f
C908 porb.t2 dvss 0.018111f
C909 porb.t5 dvss 0.018111f
C910 porb.n12 dvss 0.040174f
C911 porb.t19 dvss 0.025356f
C912 porb.t24 dvss 0.025356f
C913 porb.n13 dvss 0.0528f
C914 porb.t37 dvss 0.025356f
C915 porb.t41 dvss 0.025356f
C916 porb.n14 dvss 0.052529f
C917 porb.n15 dvss 0.52367f
C918 porb.t13 dvss 0.018111f
C919 porb.t9 dvss 0.018111f
C920 porb.n16 dvss 0.040174f
C921 porb.t46 dvss 0.025356f
C922 porb.t32 dvss 0.025356f
C923 porb.n17 dvss 0.0528f
C924 porb.t31 dvss 0.025356f
C925 porb.t17 dvss 0.025356f
C926 porb.n18 dvss 0.052529f
C927 porb.n19 dvss 0.52367f
C928 porb.t1 dvss 0.018111f
C929 porb.t12 dvss 0.018111f
C930 porb.n20 dvss 0.040174f
C931 porb.t18 dvss 0.025356f
C932 porb.t40 dvss 0.025356f
C933 porb.n21 dvss 0.0528f
C934 porb.t36 dvss 0.025356f
C935 porb.t26 dvss 0.025356f
C936 porb.n22 dvss 0.052529f
C937 porb.n23 dvss 0.52367f
C938 porb.t6 dvss 0.018111f
C939 porb.t15 dvss 0.018111f
C940 porb.n24 dvss 0.040174f
C941 porb.t27 dvss 0.025356f
C942 porb.t34 dvss 0.025356f
C943 porb.n25 dvss 0.0528f
C944 porb.t44 dvss 0.025356f
C945 porb.t20 dvss 0.025356f
C946 porb.n26 dvss 0.052529f
C947 porb.n27 dvss 0.52367f
C948 porb.t3 dvss 0.018111f
C949 porb.t11 dvss 0.018111f
C950 porb.n28 dvss 0.040174f
C951 porb.t22 dvss 0.025356f
C952 porb.t39 dvss 0.025356f
C953 porb.n29 dvss 0.0528f
C954 porb.t38 dvss 0.025356f
C955 porb.t23 dvss 0.025356f
C956 porb.n30 dvss 0.052529f
C957 porb.n31 dvss 0.52367f
C958 porb.n32 dvss 0.56314f
C959 porb.n33 dvss 0.624258f
C960 porb.n34 dvss 0.624258f
C961 porb.n35 dvss 0.624258f
C962 porb.n36 dvss 0.624258f
C963 porb.n37 dvss 0.624258f
C964 porb.n38 dvss 0.622292f
C965 porb.n39 dvss 0.656756f
C966 a_35469_n289052.n0 dvss 1.8989f
C967 a_35469_n289052.n1 dvss 1.889f
C968 a_35469_n289052.t14 dvss 0.021433f
C969 a_35469_n289052.t23 dvss 0.015309f
C970 a_35469_n289052.t15 dvss 0.015309f
C971 a_35469_n289052.n2 dvss 0.033959f
C972 a_35469_n289052.t16 dvss 0.015309f
C973 a_35469_n289052.t7 dvss 0.015309f
C974 a_35469_n289052.n3 dvss 0.033959f
C975 a_35469_n289052.t18 dvss 0.021433f
C976 a_35469_n289052.t10 dvss 0.021433f
C977 a_35469_n289052.n4 dvss 0.044631f
C978 a_35469_n289052.t8 dvss 0.021433f
C979 a_35469_n289052.t1 dvss 0.021433f
C980 a_35469_n289052.n5 dvss 0.044402f
C981 a_35469_n289052.t5 dvss 0.015309f
C982 a_35469_n289052.t9 dvss 0.015309f
C983 a_35469_n289052.n6 dvss 0.033959f
C984 a_35469_n289052.t4 dvss 0.021433f
C985 a_35469_n289052.t3 dvss 0.021433f
C986 a_35469_n289052.n7 dvss 0.044631f
C987 a_35469_n289052.t22 dvss 0.021433f
C988 a_35469_n289052.t19 dvss 0.021433f
C989 a_35469_n289052.n8 dvss 0.044402f
C990 a_35469_n289052.t13 dvss 0.015309f
C991 a_35469_n289052.t11 dvss 0.015309f
C992 a_35469_n289052.n9 dvss 0.033959f
C993 a_35469_n289052.t17 dvss 0.021433f
C994 a_35469_n289052.t20 dvss 0.021433f
C995 a_35469_n289052.n10 dvss 0.044631f
C996 a_35469_n289052.t21 dvss 0.021433f
C997 a_35469_n289052.t12 dvss 0.021433f
C998 a_35469_n289052.n11 dvss 0.044402f
C999 a_35469_n289052.t54 dvss 0.016701f
C1000 a_35469_n289052.t62 dvss 0.016701f
C1001 a_35469_n289052.t47 dvss 0.016701f
C1002 a_35469_n289052.t27 dvss 0.016701f
C1003 a_35469_n289052.t59 dvss 0.016701f
C1004 a_35469_n289052.t38 dvss 0.016701f
C1005 a_35469_n289052.t66 dvss 0.016701f
C1006 a_35469_n289052.t49 dvss 0.035041f
C1007 a_35469_n289052.n12 dvss 0.099069f
C1008 a_35469_n289052.n13 dvss 0.068808f
C1009 a_35469_n289052.n14 dvss 0.068808f
C1010 a_35469_n289052.n15 dvss 0.068808f
C1011 a_35469_n289052.n16 dvss 0.068808f
C1012 a_35469_n289052.n17 dvss 0.068808f
C1013 a_35469_n289052.n18 dvss 0.054111f
C1014 a_35469_n289052.t28 dvss 0.016701f
C1015 a_35469_n289052.t43 dvss 0.016701f
C1016 a_35469_n289052.t63 dvss 0.016701f
C1017 a_35469_n289052.t32 dvss 0.016701f
C1018 a_35469_n289052.t51 dvss 0.016701f
C1019 a_35469_n289052.t24 dvss 0.016701f
C1020 a_35469_n289052.t61 dvss 0.016701f
C1021 a_35469_n289052.t34 dvss 0.035041f
C1022 a_35469_n289052.n19 dvss 0.099069f
C1023 a_35469_n289052.n20 dvss 0.068808f
C1024 a_35469_n289052.n21 dvss 0.068808f
C1025 a_35469_n289052.n22 dvss 0.068808f
C1026 a_35469_n289052.n23 dvss 0.068808f
C1027 a_35469_n289052.n24 dvss 0.068808f
C1028 a_35469_n289052.n25 dvss 0.054111f
C1029 a_35469_n289052.n26 dvss 0.289399f
C1030 a_35469_n289052.t58 dvss 0.041474f
C1031 a_35469_n289052.t35 dvss 0.044675f
C1032 a_35469_n289052.t68 dvss 0.041474f
C1033 a_35469_n289052.t40 dvss 0.044675f
C1034 a_35469_n289052.t50 dvss 0.041474f
C1035 a_35469_n289052.t25 dvss 0.044675f
C1036 a_35469_n289052.t31 dvss 0.041474f
C1037 a_35469_n289052.t52 dvss 0.044675f
C1038 a_35469_n289052.t57 dvss 0.041474f
C1039 a_35469_n289052.t33 dvss 0.044675f
C1040 a_35469_n289052.t42 dvss 0.041474f
C1041 a_35469_n289052.t65 dvss 0.044675f
C1042 a_35469_n289052.t71 dvss 0.041474f
C1043 a_35469_n289052.t45 dvss 0.044675f
C1044 a_35469_n289052.t53 dvss 0.041474f
C1045 a_35469_n289052.t29 dvss 0.060555f
C1046 a_35469_n289052.n27 dvss 0.1096f
C1047 a_35469_n289052.n28 dvss 0.072844f
C1048 a_35469_n289052.n29 dvss 0.072844f
C1049 a_35469_n289052.n30 dvss 0.072844f
C1050 a_35469_n289052.n31 dvss 0.072844f
C1051 a_35469_n289052.n32 dvss 0.072844f
C1052 a_35469_n289052.n33 dvss 0.058147f
C1053 a_35469_n289052.t26 dvss 0.041474f
C1054 a_35469_n289052.t48 dvss 0.044675f
C1055 a_35469_n289052.t46 dvss 0.041474f
C1056 a_35469_n289052.t70 dvss 0.044675f
C1057 a_35469_n289052.t69 dvss 0.041474f
C1058 a_35469_n289052.t41 dvss 0.044675f
C1059 a_35469_n289052.t36 dvss 0.041474f
C1060 a_35469_n289052.t56 dvss 0.044675f
C1061 a_35469_n289052.t55 dvss 0.041474f
C1062 a_35469_n289052.t30 dvss 0.044675f
C1063 a_35469_n289052.t44 dvss 0.041474f
C1064 a_35469_n289052.t67 dvss 0.044675f
C1065 a_35469_n289052.t64 dvss 0.041474f
C1066 a_35469_n289052.t39 dvss 0.044675f
C1067 a_35469_n289052.t37 dvss 0.041474f
C1068 a_35469_n289052.t60 dvss 0.060555f
C1069 a_35469_n289052.n34 dvss 0.1096f
C1070 a_35469_n289052.n35 dvss 0.072844f
C1071 a_35469_n289052.n36 dvss 0.072844f
C1072 a_35469_n289052.n37 dvss 0.072844f
C1073 a_35469_n289052.n38 dvss 0.072844f
C1074 a_35469_n289052.n39 dvss 0.072844f
C1075 a_35469_n289052.n40 dvss 0.058147f
C1076 a_35469_n289052.n41 dvss 0.284893f
C1077 a_35469_n289052.n42 dvss 1.908f
C1078 a_35469_n289052.t6 dvss 0.021433f
C1079 a_35469_n289052.t2 dvss 0.021433f
C1080 a_35469_n289052.n43 dvss 0.044402f
C1081 a_35469_n289052.n44 dvss 0.044631f
C1082 a_35469_n289052.t0 dvss 0.021433f
C1083 x1.vo.t3 dvss 0.052804f
C1084 x1.vo.t4 dvss 0.10768f
C1085 x1.vo.n0 dvss 0.230099f
C1086 x1.vo.t5 dvss 12.3449f
C1087 x1.vo.n1 dvss 0.135637f
C1088 x1.vo.t2 dvss 0.070554f
C1089 x1.vo.t1 dvss 0.034431f
C1090 x1.vo.t0 dvss 0.032156f
C1091 x1.vo.n2 dvss 0.243288f
C1092 x1.vo.n3 dvss 0.248455f
C1093 x1.vt.t3 dvss 0.263269f
C1094 x1.vt.t2 dvss 0.164219f
C1095 x1.vt.t0 dvss 0.219002f
C1096 x1.vt.n0 dvss 0.892457f
C1097 x1.vt.t1 dvss 19.7699f
C1098 a_28094_n290278.t4 dvss 0.022694f
C1099 a_28094_n290278.t2 dvss 0.022694f
C1100 a_28094_n290278.t5 dvss 0.022694f
C1101 a_28094_n290278.n0 dvss 0.047876f
C1102 a_28094_n290278.t9 dvss 0.086108f
C1103 a_28094_n290278.t8 dvss 0.084311f
C1104 a_28094_n290278.n1 dvss 1.22225f
C1105 a_28094_n290278.n2 dvss 0.886586f
C1106 a_28094_n290278.t3 dvss 0.022694f
C1107 a_28094_n290278.t6 dvss 0.022694f
C1108 a_28094_n290278.n3 dvss 0.047893f
C1109 a_28094_n290278.t0 dvss 0.022694f
C1110 a_28094_n290278.t1 dvss 0.022694f
C1111 a_28094_n290278.n4 dvss 0.049537f
C1112 a_28094_n290278.n5 dvss 1.16932f
C1113 a_28094_n290278.n6 dvss 0.676718f
C1114 a_28094_n290278.n7 dvss 0.047855f
C1115 a_28094_n290278.t7 dvss 0.022694f
C1116 x2.vbp1.n0 dvss 0.349388f
C1117 x2.vbp1.n1 dvss 1.25652f
C1118 x2.vbp1.t30 dvss 60.755898f
C1119 x2.vbp1.t8 dvss 0.07584f
C1120 x2.vbp1.t36 dvss 0.074618f
C1121 x2.vbp1.n2 dvss 0.143216f
C1122 x2.vbp1.t10 dvss 0.07584f
C1123 x2.vbp1.t35 dvss 0.074618f
C1124 x2.vbp1.n3 dvss 0.143216f
C1125 x2.vbp1.t18 dvss 0.07584f
C1126 x2.vbp1.t32 dvss 0.074618f
C1127 x2.vbp1.n4 dvss 0.143216f
C1128 x2.vbp1.t12 dvss 0.07584f
C1129 x2.vbp1.t34 dvss 0.074618f
C1130 x2.vbp1.n5 dvss 0.14268f
C1131 x2.vbp1.t6 dvss 0.07584f
C1132 x2.vbp1.t37 dvss 0.074618f
C1133 x2.vbp1.n6 dvss 0.14268f
C1134 x2.vbp1.t31 dvss 0.074982f
C1135 x2.vbp1.t39 dvss 0.075403f
C1136 x2.vbp1.n7 dvss 0.172631f
C1137 x2.vbp1.t28 dvss 0.025125f
C1138 x2.vbp1.t29 dvss 0.025434f
C1139 x2.vbp1.n8 dvss 0.302615f
C1140 x2.vbp1.n9 dvss 0.014306f
C1141 x2.vbp1.n10 dvss 0.014226f
C1142 x2.vbp1.n11 dvss 0.014636f
C1143 x2.vbp1.n12 dvss 0.45365f
C1144 x2.vbp1.n13 dvss 0.014147f
C1145 x2.vbp1.n14 dvss 0.01415f
C1146 x2.vbp1.n15 dvss 0.140448f
C1147 x2.vbp1.n16 dvss 0.01415f
C1148 x2.vbp1.n17 dvss 0.140224f
C1149 x2.vbp1.n18 dvss 0.01415f
C1150 x2.vbp1.n19 dvss 0.123921f
C1151 x2.vbp1.n20 dvss 0.056882f
C1152 x2.vbp1.n21 dvss 0.062153f
C1153 x2.vbp1.n22 dvss 0.04547f
C1154 x2.vbp1.n23 dvss 0.045271f
C1155 x2.vbp1.n24 dvss 0.045293f
C1156 x2.vbp1.n25 dvss 0.043166f
C1157 x2.vbp1.t14 dvss 0.07584f
C1158 x2.vbp1.t33 dvss 0.074618f
C1159 x2.vbp1.n26 dvss 0.143216f
C1160 x2.vbp1.t20 dvss 0.07584f
C1161 x2.vbp1.t40 dvss 0.074618f
C1162 x2.vbp1.n27 dvss 0.143216f
C1163 x2.vbp1.t4 dvss 0.07584f
C1164 x2.vbp1.t38 dvss 0.074618f
C1165 x2.vbp1.n28 dvss 0.143216f
C1166 x2.vbp1.t24 dvss 0.07584f
C1167 x2.vbp1.t2 dvss 0.074618f
C1168 x2.vbp1.n29 dvss 0.143216f
C1169 x2.vbp1.t16 dvss 0.07584f
C1170 x2.vbp1.t22 dvss 0.074618f
C1171 x2.vbp1.n30 dvss 0.143216f
C1172 x2.vbp1.t0 dvss 0.075296f
C1173 x2.vbp1.t26 dvss 0.075773f
C1174 x2.vbp1.n31 dvss 0.196362f
C1175 x2.vbp1.n32 dvss 0.045363f
C1176 x2.vbp1.n33 dvss 0.045184f
C1177 x2.vbp1.n34 dvss 0.045328f
C1178 x2.vbp1.n35 dvss 0.045219f
C1179 por.t36 dvss 0.019758f
C1180 por.t23 dvss 0.019758f
C1181 por.n0 dvss 0.041144f
C1182 por.t44 dvss 0.019758f
C1183 por.t30 dvss 0.019758f
C1184 por.n1 dvss 0.040933f
C1185 por.n2 dvss 0.406695f
C1186 por.t1 dvss 0.014113f
C1187 por.t10 dvss 0.014113f
C1188 por.n3 dvss 0.031265f
C1189 por.t45 dvss 0.019758f
C1190 por.t31 dvss 0.019758f
C1191 por.n4 dvss 0.041144f
C1192 por.t19 dvss 0.019758f
C1193 por.t38 dvss 0.019758f
C1194 por.n5 dvss 0.040933f
C1195 por.n6 dvss 0.408064f
C1196 por.t5 dvss 0.014113f
C1197 por.t14 dvss 0.014113f
C1198 por.n7 dvss 0.031305f
C1199 por.t20 dvss 0.019758f
C1200 por.t39 dvss 0.019758f
C1201 por.n8 dvss 0.041144f
C1202 por.t27 dvss 0.019758f
C1203 por.t47 dvss 0.019758f
C1204 por.n9 dvss 0.040933f
C1205 por.n10 dvss 0.408064f
C1206 por.t7 dvss 0.014113f
C1207 por.t3 dvss 0.014113f
C1208 por.n11 dvss 0.031305f
C1209 por.t24 dvss 0.019758f
C1210 por.t33 dvss 0.019758f
C1211 por.n12 dvss 0.041144f
C1212 por.t32 dvss 0.019758f
C1213 por.t40 dvss 0.019758f
C1214 por.n13 dvss 0.040933f
C1215 por.n14 dvss 0.408064f
C1216 por.t11 dvss 0.014113f
C1217 por.t15 dvss 0.014113f
C1218 por.n15 dvss 0.031305f
C1219 por.t18 dvss 0.019758f
C1220 por.t41 dvss 0.019758f
C1221 por.n16 dvss 0.041144f
C1222 por.t25 dvss 0.019758f
C1223 por.t16 dvss 0.019758f
C1224 por.n17 dvss 0.040933f
C1225 por.n18 dvss 0.408064f
C1226 por.t8 dvss 0.014113f
C1227 por.t2 dvss 0.014113f
C1228 por.n19 dvss 0.031305f
C1229 por.t26 dvss 0.019758f
C1230 por.t46 dvss 0.019758f
C1231 por.n20 dvss 0.041144f
C1232 por.t34 dvss 0.019758f
C1233 por.t21 dvss 0.019758f
C1234 por.n21 dvss 0.040933f
C1235 por.n22 dvss 0.408064f
C1236 por.t12 dvss 0.014113f
C1237 por.t6 dvss 0.014113f
C1238 por.n23 dvss 0.031305f
C1239 por.t35 dvss 0.019758f
C1240 por.t22 dvss 0.019758f
C1241 por.n24 dvss 0.041144f
C1242 por.t42 dvss 0.019758f
C1243 por.t28 dvss 0.019758f
C1244 por.n25 dvss 0.040933f
C1245 por.n26 dvss 0.408064f
C1246 por.t0 dvss 0.014113f
C1247 por.t9 dvss 0.014113f
C1248 por.n27 dvss 0.031305f
C1249 por.t43 dvss 0.019758f
C1250 por.t29 dvss 0.019758f
C1251 por.n28 dvss 0.041144f
C1252 por.t17 dvss 0.019758f
C1253 por.t37 dvss 0.019758f
C1254 por.n29 dvss 0.040933f
C1255 por.n30 dvss 0.408064f
C1256 por.t4 dvss 0.014113f
C1257 por.t13 dvss 0.014113f
C1258 por.n31 dvss 0.031305f
C1259 por.n32 dvss 0.438821f
C1260 por.n33 dvss 0.486446f
C1261 por.n34 dvss 0.486446f
C1262 por.n35 dvss 0.486446f
C1263 por.n36 dvss 0.486446f
C1264 por.n37 dvss 0.486446f
C1265 por.n38 dvss 0.484914f
C1266 por.n39 dvss 0.48569f
C1267 por.n40 dvss 0.858126f
C1268 a_35454_n291454.n0 dvss 0.438871f
C1269 a_35454_n291454.t17 dvss 0.018705f
C1270 a_35454_n291454.t1 dvss 0.013361f
C1271 a_35454_n291454.t7 dvss 0.013361f
C1272 a_35454_n291454.n1 dvss 0.029637f
C1273 a_35454_n291454.t20 dvss 0.018705f
C1274 a_35454_n291454.t11 dvss 0.018705f
C1275 a_35454_n291454.n2 dvss 0.038951f
C1276 a_35454_n291454.t22 dvss 0.018705f
C1277 a_35454_n291454.t16 dvss 0.018705f
C1278 a_35454_n291454.n3 dvss 0.038751f
C1279 a_35454_n291454.n4 dvss 0.386315f
C1280 a_35454_n291454.t0 dvss 0.013361f
C1281 a_35454_n291454.t4 dvss 0.013361f
C1282 a_35454_n291454.n5 dvss 0.029637f
C1283 a_35454_n291454.t15 dvss 0.018705f
C1284 a_35454_n291454.t9 dvss 0.018705f
C1285 a_35454_n291454.n6 dvss 0.038951f
C1286 a_35454_n291454.t19 dvss 0.018705f
C1287 a_35454_n291454.t14 dvss 0.018705f
C1288 a_35454_n291454.n7 dvss 0.038751f
C1289 a_35454_n291454.n8 dvss 0.386315f
C1290 a_35454_n291454.t6 dvss 0.013361f
C1291 a_35454_n291454.t2 dvss 0.013361f
C1292 a_35454_n291454.n9 dvss 0.029637f
C1293 a_35454_n291454.t8 dvss 0.018705f
C1294 a_35454_n291454.t13 dvss 0.018705f
C1295 a_35454_n291454.n10 dvss 0.038951f
C1296 a_35454_n291454.t12 dvss 0.018705f
C1297 a_35454_n291454.t18 dvss 0.018705f
C1298 a_35454_n291454.n11 dvss 0.038751f
C1299 a_35454_n291454.n12 dvss 0.386315f
C1300 a_35454_n291454.t3 dvss 0.013361f
C1301 a_35454_n291454.t5 dvss 0.013361f
C1302 a_35454_n291454.n13 dvss 0.029637f
C1303 a_35454_n291454.t44 dvss 0.036196f
C1304 a_35454_n291454.t34 dvss 0.038989f
C1305 a_35454_n291454.t57 dvss 0.036196f
C1306 a_35454_n291454.t46 dvss 0.038989f
C1307 a_35454_n291454.t36 dvss 0.036196f
C1308 a_35454_n291454.t24 dvss 0.038989f
C1309 a_35454_n291454.t62 dvss 0.036196f
C1310 a_35454_n291454.t53 dvss 0.038989f
C1311 a_35454_n291454.t48 dvss 0.036196f
C1312 a_35454_n291454.t37 dvss 0.038989f
C1313 a_35454_n291454.t27 dvss 0.036196f
C1314 a_35454_n291454.t63 dvss 0.038989f
C1315 a_35454_n291454.t59 dvss 0.036196f
C1316 a_35454_n291454.t49 dvss 0.038989f
C1317 a_35454_n291454.t39 dvss 0.036196f
C1318 a_35454_n291454.t28 dvss 0.052848f
C1319 a_35454_n291454.n14 dvss 0.095651f
C1320 a_35454_n291454.n15 dvss 0.063573f
C1321 a_35454_n291454.n16 dvss 0.063573f
C1322 a_35454_n291454.n17 dvss 0.063573f
C1323 a_35454_n291454.n18 dvss 0.063573f
C1324 a_35454_n291454.n19 dvss 0.063573f
C1325 a_35454_n291454.n20 dvss 0.050747f
C1326 a_35454_n291454.t64 dvss 0.036196f
C1327 a_35454_n291454.t55 dvss 0.038989f
C1328 a_35454_n291454.t32 dvss 0.036196f
C1329 a_35454_n291454.t69 dvss 0.038989f
C1330 a_35454_n291454.t54 dvss 0.036196f
C1331 a_35454_n291454.t42 dvss 0.038989f
C1332 a_35454_n291454.t25 dvss 0.036196f
C1333 a_35454_n291454.t61 dvss 0.038989f
C1334 a_35454_n291454.t41 dvss 0.036196f
C1335 a_35454_n291454.t30 dvss 0.038989f
C1336 a_35454_n291454.t60 dvss 0.036196f
C1337 a_35454_n291454.t51 dvss 0.038989f
C1338 a_35454_n291454.t29 dvss 0.036196f
C1339 a_35454_n291454.t66 dvss 0.038989f
C1340 a_35454_n291454.t50 dvss 0.036196f
C1341 a_35454_n291454.t38 dvss 0.052848f
C1342 a_35454_n291454.n21 dvss 0.095651f
C1343 a_35454_n291454.n22 dvss 0.063573f
C1344 a_35454_n291454.n23 dvss 0.063573f
C1345 a_35454_n291454.n24 dvss 0.063573f
C1346 a_35454_n291454.n25 dvss 0.063573f
C1347 a_35454_n291454.n26 dvss 0.063573f
C1348 a_35454_n291454.n27 dvss 0.050747f
C1349 a_35454_n291454.n28 dvss 0.248634f
C1350 a_35454_n291454.t26 dvss 0.014575f
C1351 a_35454_n291454.t40 dvss 0.014575f
C1352 a_35454_n291454.t67 dvss 0.014575f
C1353 a_35454_n291454.t52 dvss 0.014575f
C1354 a_35454_n291454.t31 dvss 0.014575f
C1355 a_35454_n291454.t58 dvss 0.014575f
C1356 a_35454_n291454.t43 dvss 0.014575f
C1357 a_35454_n291454.t70 dvss 0.030581f
C1358 a_35454_n291454.n29 dvss 0.08646f
C1359 a_35454_n291454.n30 dvss 0.060051f
C1360 a_35454_n291454.n31 dvss 0.060051f
C1361 a_35454_n291454.n32 dvss 0.060051f
C1362 a_35454_n291454.n33 dvss 0.060051f
C1363 a_35454_n291454.n34 dvss 0.060051f
C1364 a_35454_n291454.n35 dvss 0.047224f
C1365 a_35454_n291454.t47 dvss 0.014575f
C1366 a_35454_n291454.t68 dvss 0.014575f
C1367 a_35454_n291454.t35 dvss 0.014575f
C1368 a_35454_n291454.t56 dvss 0.014575f
C1369 a_35454_n291454.t71 dvss 0.014575f
C1370 a_35454_n291454.t45 dvss 0.014575f
C1371 a_35454_n291454.t65 dvss 0.014575f
C1372 a_35454_n291454.t33 dvss 0.030581f
C1373 a_35454_n291454.n36 dvss 0.08646f
C1374 a_35454_n291454.n37 dvss 0.060051f
C1375 a_35454_n291454.n38 dvss 0.060051f
C1376 a_35454_n291454.n39 dvss 0.060051f
C1377 a_35454_n291454.n40 dvss 0.060051f
C1378 a_35454_n291454.n41 dvss 0.060051f
C1379 a_35454_n291454.n42 dvss 0.047224f
C1380 a_35454_n291454.n43 dvss 0.252567f
C1381 a_35454_n291454.n44 dvss 1.66517f
C1382 a_35454_n291454.n45 dvss 0.445725f
C1383 a_35454_n291454.n46 dvss 0.460519f
C1384 a_35454_n291454.n47 dvss 0.415432f
C1385 a_35454_n291454.t10 dvss 0.018705f
C1386 a_35454_n291454.t21 dvss 0.018705f
C1387 a_35454_n291454.n48 dvss 0.038751f
C1388 a_35454_n291454.n49 dvss 0.386315f
C1389 a_35454_n291454.n50 dvss 0.038951f
C1390 a_35454_n291454.t23 dvss 0.018705f
C1391 a_34073_n287091.n0 dvss 0.283068f
C1392 a_34073_n287091.n1 dvss 1.09949f
C1393 a_34073_n287091.n2 dvss 0.064289f
C1394 a_34073_n287091.n3 dvss 0.196887f
C1395 a_34073_n287091.n4 dvss 0.374447f
C1396 a_34073_n287091.t1 dvss 0.097396f
C1397 a_34073_n287091.t2 dvss 0.058657f
C1398 a_34073_n287091.t0 dvss 0.097211f
C1399 a_34073_n287091.t5 dvss 0.168419f
C1400 a_34073_n287091.t9 dvss 0.168259f
C1401 a_34073_n287091.t8 dvss 0.125353f
C1402 a_34073_n287091.t4 dvss 1.56507f
C1403 a_34073_n287091.n5 dvss 0.329321f
C1404 a_34073_n287091.t7 dvss 0.167622f
C1405 a_34073_n287091.n6 dvss 0.178025f
C1406 a_34073_n287091.t6 dvss 0.167695f
C1407 a_34073_n287091.t3 dvss 0.058796f
C1408 porb_h[1].t9 dvss 0.015201f
C1409 porb_h[1].t6 dvss 0.015201f
C1410 porb_h[1].n0 dvss 0.062532f
C1411 porb_h[1].t21 dvss 0.030403f
C1412 porb_h[1].t20 dvss 0.030403f
C1413 porb_h[1].n1 dvss 0.072126f
C1414 porb_h[1].n2 dvss 0.231154f
C1415 porb_h[1].n3 dvss 0.017882f
C1416 porb_h[1].n4 dvss 0.018365f
C1417 porb_h[1].n5 dvss 0.133518f
C1418 porb_h[1].t0 dvss 0.015201f
C1419 porb_h[1].t15 dvss 0.015201f
C1420 porb_h[1].n6 dvss 0.062532f
C1421 porb_h[1].t29 dvss 0.030403f
C1422 porb_h[1].t28 dvss 0.030403f
C1423 porb_h[1].n7 dvss 0.072126f
C1424 porb_h[1].n8 dvss 0.231154f
C1425 porb_h[1].n9 dvss 0.208129f
C1426 porb_h[1].t11 dvss 0.015201f
C1427 porb_h[1].t5 dvss 0.015201f
C1428 porb_h[1].n10 dvss 0.062532f
C1429 porb_h[1].t25 dvss 0.030403f
C1430 porb_h[1].t17 dvss 0.030403f
C1431 porb_h[1].n11 dvss 0.072126f
C1432 porb_h[1].n12 dvss 0.231154f
C1433 porb_h[1].n13 dvss 0.238329f
C1434 porb_h[1].t12 dvss 0.015201f
C1435 porb_h[1].t4 dvss 0.015201f
C1436 porb_h[1].n14 dvss 0.062532f
C1437 porb_h[1].t24 dvss 0.030403f
C1438 porb_h[1].t16 dvss 0.030403f
C1439 porb_h[1].n15 dvss 0.072126f
C1440 porb_h[1].n16 dvss 0.231154f
C1441 porb_h[1].n17 dvss 0.238329f
C1442 porb_h[1].t7 dvss 0.015201f
C1443 porb_h[1].t13 dvss 0.015201f
C1444 porb_h[1].n18 dvss 0.062532f
C1445 porb_h[1].t19 dvss 0.030403f
C1446 porb_h[1].t26 dvss 0.030403f
C1447 porb_h[1].n19 dvss 0.072126f
C1448 porb_h[1].n20 dvss 0.231154f
C1449 porb_h[1].n21 dvss 0.238329f
C1450 porb_h[1].t14 dvss 0.015201f
C1451 porb_h[1].t8 dvss 0.015201f
C1452 porb_h[1].n22 dvss 0.062532f
C1453 porb_h[1].t27 dvss 0.030403f
C1454 porb_h[1].t22 dvss 0.030403f
C1455 porb_h[1].n23 dvss 0.072126f
C1456 porb_h[1].n24 dvss 0.231154f
C1457 porb_h[1].n25 dvss 0.238329f
C1458 porb_h[1].t10 dvss 0.015201f
C1459 porb_h[1].t2 dvss 0.015201f
C1460 porb_h[1].n26 dvss 0.062532f
C1461 porb_h[1].t23 dvss 0.030403f
C1462 porb_h[1].t31 dvss 0.030403f
C1463 porb_h[1].n27 dvss 0.072126f
C1464 porb_h[1].n28 dvss 0.231154f
C1465 porb_h[1].n29 dvss 0.238329f
C1466 porb_h[1].t3 dvss 0.015201f
C1467 porb_h[1].t1 dvss 0.015201f
C1468 porb_h[1].n30 dvss 0.062532f
C1469 porb_h[1].t18 dvss 0.030403f
C1470 porb_h[1].t30 dvss 0.030403f
C1471 porb_h[1].n31 dvss 0.072126f
C1472 porb_h[1].n32 dvss 0.231154f
C1473 porb_h[1].n33 dvss 0.467605f
C1474 porb_h[1].n34 dvss 0.262666f
C1475 porb_h[1].n35 dvss 0.802488f
C1476 a_25567_n288267.n0 dvss 0.034229f
C1477 a_25567_n288267.n1 dvss 0.129336f
C1478 a_25567_n288267.t0 dvss 3.42214f
C1479 a_25251_n288267.n0 dvss 0.050875f
C1480 a_25251_n288267.n1 dvss 0.023453f
C1481 a_25251_n288267.n2 dvss 0.030698f
C1482 a_25251_n288267.t0 dvss 3.08131f
C1483 avdd.t15 dvss 0.030711f
C1484 avdd.n0 dvss 0.034562f
C1485 avdd.n1 dvss 0.018569f
C1486 avdd.n2 dvss 0.029051f
C1487 avdd.n3 dvss 0.033042f
C1488 avdd.n4 dvss 0.312029f
C1489 avdd.n5 dvss 0.301913f
C1490 avdd.n6 dvss 0.03085f
C1491 avdd.n7 dvss 0.033042f
C1492 avdd.n8 dvss 0.01966f
C1493 avdd.n9 dvss 0.033042f
C1494 avdd.n10 dvss 0.301913f
C1495 avdd.n11 dvss 0.03085f
C1496 avdd.n13 dvss 0.020191f
C1497 avdd.t14 dvss 0.325707f
C1498 avdd.n14 dvss 0.034568f
C1499 avdd.n15 dvss 0.312029f
C1500 avdd.n16 dvss 0.028122f
C1501 avdd.n17 dvss 0.018569f
C1502 avdd.n18 dvss 0.062388f
C1503 avdd.n19 dvss 0.090858f
C1504 avdd.n20 dvss 0.034568f
C1505 avdd.n21 dvss 0.033042f
C1506 avdd.n22 dvss 0.017617f
C1507 avdd.t8 dvss 0.301913f
C1508 avdd.n23 dvss 0.017617f
C1509 avdd.n24 dvss 0.010327f
C1510 avdd.n25 dvss 0.01966f
C1511 avdd.n26 dvss 0.020191f
C1512 avdd.n27 dvss 0.034568f
C1513 avdd.t13 dvss 0.325707f
C1514 avdd.n29 dvss 0.034568f
C1515 avdd.n30 dvss 0.099412f
C1516 avdd.n31 dvss 0.054403f
C1517 avdd.n32 dvss 0.039918f
C1518 avdd.n33 dvss 0.038743f
C1519 avdd.t95 dvss 0.060449f
C1520 avdd.n34 dvss 0.111445f
C1521 avdd.t10 dvss 0.060449f
C1522 avdd.n35 dvss 0.216601f
C1523 avdd.n36 dvss 0.154939f
C1524 avdd.t112 dvss 0.060449f
C1525 avdd.n37 dvss 0.030809f
C1526 avdd.n38 dvss 0.041312f
C1527 avdd.n39 dvss 0.041312f
C1528 avdd.n40 dvss 0.423408f
C1529 avdd.n41 dvss 0.017617f
C1530 avdd.n42 dvss 0.041312f
C1531 avdd.n43 dvss 0.16754f
C1532 avdd.n44 dvss 0.066308f
C1533 avdd.n45 dvss 0.399719f
C1534 avdd.n46 dvss 0.047391f
C1535 avdd.n47 dvss 0.041312f
C1536 avdd.n48 dvss 0.06281f
C1537 avdd.n49 dvss 0.054586f
C1538 avdd.n50 dvss 0.054586f
C1539 avdd.n51 dvss 0.274658f
C1540 avdd.n52 dvss 0.320459f
C1541 avdd.n53 dvss 0.220376f
C1542 avdd.t24 dvss 0.014999f
C1543 avdd.n55 dvss 0.023318f
C1544 avdd.n56 dvss 0.019241f
C1545 avdd.n57 dvss 0.049047f
C1546 avdd.n58 dvss 0.049047f
C1547 avdd.n59 dvss 0.133125f
C1548 avdd.t12 dvss 0.014999f
C1549 avdd.t19 dvss 0.014632f
C1550 avdd.n60 dvss 0.032418f
C1551 avdd.t17 dvss 0.01474f
C1552 avdd.t16 dvss 0.07814f
C1553 avdd.n61 dvss 0.104197f
C1554 avdd.n62 dvss 0.060643f
C1555 avdd.t18 dvss 0.078058f
C1556 avdd.n63 dvss 0.069419f
C1557 avdd.n64 dvss 0.080055f
C1558 avdd.t27 dvss 0.029997f
C1559 avdd.n65 dvss 0.052166f
C1560 avdd.n66 dvss 0.314266f
C1561 avdd.n67 dvss 0.251809f
C1562 avdd.n68 dvss 0.410116f
C1563 avdd.n69 dvss 0.017362f
C1564 avdd.n70 dvss 0.018142f
C1565 avdd.n71 dvss 0.067585f
C1566 avdd.n72 dvss 0.01722f
C1567 avdd.n73 dvss 0.255918f
C1568 avdd.t11 dvss 0.186743f
C1569 avdd.n74 dvss 0.089447f
C1570 avdd.t23 dvss 0.165306f
C1571 avdd.n75 dvss 0.196412f
C1572 avdd.n76 dvss 0.049209f
C1573 avdd.n77 dvss 0.018258f
C1574 avdd.n78 dvss 0.056682f
C1575 avdd.n79 dvss 0.199837f
C1576 avdd.n80 dvss 0.123547f
C1577 avdd.n81 dvss 0.15619f
C1578 avdd.n82 dvss 0.055415f
C1579 avdd.t26 dvss 0.372785f
C1580 avdd.n83 dvss 0.055415f
C1581 avdd.n84 dvss 0.018615f
C1582 avdd.n85 dvss 0.046835f
C1583 avdd.n86 dvss 0.222386f
C1584 avdd.n87 dvss 0.010327f
C1585 avdd.n88 dvss 0.031028f
C1586 avdd.n89 dvss 0.025027f
C1587 avdd.n90 dvss 0.043061f
C1588 avdd.t94 dvss 0.423408f
C1589 avdd.n91 dvss 0.043061f
C1590 avdd.n92 dvss 0.13586f
C1591 avdd.n93 dvss 0.154644f
C1592 avdd.n94 dvss 0.093245f
C1593 avdd.n95 dvss 0.017617f
C1594 avdd.t9 dvss 0.423408f
C1595 avdd.n97 dvss 0.435488f
C1596 avdd.n98 dvss 0.043061f
C1597 avdd.n99 dvss 0.035006f
C1598 avdd.n100 dvss 0.120714f
C1599 avdd.n101 dvss 0.218532f
C1600 avdd.n102 dvss 0.043061f
C1601 avdd.t111 dvss 0.454775f
C1602 avdd.n103 dvss 0.423408f
C1603 avdd.n104 dvss 0.047391f
C1604 avdd.n105 dvss 0.216202f
C1605 avdd.t124 dvss 0.09778f
C1606 avdd.t123 dvss 0.097091f
C1607 avdd.n106 dvss 0.342351f
C1608 avdd.n107 dvss 0.617216f
C1609 avdd.n108 dvss 0.351349f
C1610 avdd.n109 dvss 0.281533f
C1611 avdd.n110 dvss 0.04115f
C1612 avdd.n111 dvss 1.04193f
C1613 avdd.n112 dvss 1.45664f
C1614 avdd.n113 dvss 2.16246f
C1615 avdd.n114 dvss 2.05578f
C1616 avdd.n115 dvss 1.78183f
C1617 avdd.n116 dvss 0.730237f
C1618 avdd.n117 dvss 1.04301f
C1619 avdd.n118 dvss 3.77692f
C1620 avdd.n119 dvss 1.80347f
C1621 avdd.n120 dvss 0.360913f
C1622 avdd.n121 dvss 1.61637f
C1623 avdd.n122 dvss 2.50139f
C1624 avdd.n123 dvss 0.469748f
C1625 avdd.n124 dvss 0.613173f
C1626 avdd.t89 dvss 0.011993f
C1627 avdd.t91 dvss 0.011993f
C1628 avdd.n125 dvss 0.025859f
C1629 avdd.t1 dvss 0.011993f
C1630 avdd.t3 dvss 0.011993f
C1631 avdd.n126 dvss 0.025841f
C1632 avdd.t81 dvss 0.011993f
C1633 avdd.t22 dvss 0.011993f
C1634 avdd.n127 dvss 0.02585f
C1635 avdd.t103 dvss 0.038699f
C1636 avdd.t105 dvss 0.038547f
C1637 avdd.n128 dvss 0.388909f
C1638 avdd.t109 dvss 0.038549f
C1639 avdd.n129 dvss 0.248965f
C1640 avdd.t107 dvss 0.038547f
C1641 avdd.n130 dvss 0.246575f
C1642 avdd.t79 dvss 0.038548f
C1643 avdd.n131 dvss 0.244152f
C1644 avdd.t115 dvss 0.038549f
C1645 avdd.n132 dvss 0.195437f
C1646 avdd.n133 dvss 0.285515f
C1647 avdd.n134 dvss 0.093365f
C1648 avdd.n135 dvss 0.029266f
C1649 avdd.n136 dvss 0.043062f
C1650 avdd.n137 dvss 0.043062f
C1651 avdd.t106 dvss 0.227765f
C1652 avdd.n138 dvss 0.041643f
C1653 avdd.n139 dvss 0.041643f
C1654 avdd.n140 dvss 0.060309f
C1655 avdd.n141 dvss 0.024702f
C1656 avdd.n142 dvss 0.041643f
C1657 avdd.t108 dvss 0.227765f
C1658 avdd.n143 dvss 0.041643f
C1659 avdd.n144 dvss 0.020751f
C1660 avdd.n145 dvss 0.175206f
C1661 avdd.n146 dvss 0.061095f
C1662 avdd.n147 dvss 0.438369f
C1663 avdd.t102 dvss 0.227765f
C1664 avdd.n148 dvss 0.062701f
C1665 avdd.n149 dvss 0.029047f
C1666 avdd.n150 dvss 0.043062f
C1667 avdd.n151 dvss 0.034985f
C1668 avdd.n152 dvss 0.332287f
C1669 avdd.t104 dvss 0.227765f
C1670 avdd.n153 dvss 0.123243f
C1671 avdd.n154 dvss 0.043062f
C1672 avdd.n155 dvss 0.09247f
C1673 avdd.n156 dvss 0.061005f
C1674 avdd.n157 dvss 0.0254f
C1675 avdd.n158 dvss 0.026096f
C1676 avdd.n159 dvss 0.024151f
C1677 avdd.n160 dvss 0.123243f
C1678 avdd.n161 dvss 0.024151f
C1679 avdd.n162 dvss 0.014157f
C1680 avdd.n163 dvss 0.024702f
C1681 avdd.n164 dvss 0.020751f
C1682 avdd.n165 dvss 0.034985f
C1683 avdd.n166 dvss 0.332287f
C1684 avdd.t78 dvss 0.227765f
C1685 avdd.n167 dvss 0.123243f
C1686 avdd.t114 dvss 0.253965f
C1687 avdd.n168 dvss 0.349241f
C1688 avdd.n169 dvss 0.064866f
C1689 avdd.n170 dvss 0.077696f
C1690 avdd.n171 dvss 0.182637f
C1691 avdd.n172 dvss 0.393422f
C1692 avdd.n173 dvss 0.530789f
C1693 avdd.n174 dvss 0.284097f
C1694 avdd.n175 dvss 0.0427f
C1695 avdd.n176 dvss 0.022642f
C1696 avdd.n177 dvss 0.037083f
C1697 avdd.n178 dvss 0.043297f
C1698 avdd.n179 dvss 0.373937f
C1699 avdd.t88 dvss 0.24442f
C1700 avdd.n180 dvss 0.043297f
C1701 avdd.n181 dvss 0.025672f
C1702 avdd.n182 dvss 0.043297f
C1703 avdd.t0 dvss 0.24442f
C1704 avdd.n183 dvss 0.038293f
C1705 avdd.n184 dvss 0.356586f
C1706 avdd.t2 dvss 0.24442f
C1707 avdd.n185 dvss 0.038293f
C1708 avdd.n186 dvss 0.373937f
C1709 avdd.n187 dvss 0.022642f
C1710 avdd.n188 dvss 0.093156f
C1711 avdd.n189 dvss 0.136099f
C1712 avdd.t80 dvss 0.272116f
C1713 avdd.n190 dvss 0.035971f
C1714 avdd.n191 dvss 0.026183f
C1715 avdd.n192 dvss 0.044768f
C1716 avdd.n193 dvss 0.356586f
C1717 avdd.t21 dvss 0.24442f
C1718 avdd.n194 dvss 0.132255f
C1719 avdd.n195 dvss 0.044768f
C1720 avdd.n196 dvss 0.043297f
C1721 avdd.n197 dvss 0.024151f
C1722 avdd.n198 dvss 0.132255f
C1723 avdd.n199 dvss 0.024151f
C1724 avdd.n200 dvss 0.014157f
C1725 avdd.n201 dvss 0.025672f
C1726 avdd.n202 dvss 0.026183f
C1727 avdd.n203 dvss 0.044768f
C1728 avdd.t90 dvss 0.272116f
C1729 avdd.n204 dvss 0.132255f
C1730 avdd.n205 dvss 0.044768f
C1731 avdd.n206 dvss 0.146224f
C1732 avdd.n207 dvss 0.09147f
C1733 avdd.n208 dvss 0.197147f
C1734 avdd.n209 dvss 0.531993f
C1735 avdd.n210 dvss 0.362262f
C1736 avdd.n211 dvss 0.105794f
C1737 avdd.t120 dvss 0.494574f
C1738 avdd.n212 dvss 0.081121f
C1739 avdd.n213 dvss 0.111129f
C1740 avdd.n214 dvss 0.013369f
C1741 avdd.n215 dvss 0.028342f
C1742 avdd.n221 dvss 0.017112f
C1743 avdd.n222 dvss 0.014552f
C1744 avdd.n223 dvss 0.077636f
C1745 avdd.n224 dvss 0.012834f
C1746 avdd.n225 dvss 0.014552f
C1747 avdd.n226 dvss 0.017112f
C1748 avdd.n230 dvss 0.014552f
C1749 avdd.n231 dvss 0.077636f
C1750 avdd.n232 dvss 0.012834f
C1751 avdd.n233 dvss 0.014552f
C1752 avdd.n234 dvss 0.022459f
C1753 avdd.t30 dvss 0.059823f
C1754 avdd.t66 dvss 0.059823f
C1755 avdd.n243 dvss 0.014552f
C1756 avdd.n244 dvss 0.077636f
C1757 avdd.n245 dvss 0.014552f
C1758 avdd.n246 dvss 0.077636f
C1759 avdd.n247 dvss 0.012834f
C1760 avdd.n248 dvss 0.014552f
C1761 avdd.n250 dvss 0.015508f
C1762 avdd.n251 dvss 0.077635f
C1763 avdd.n252 dvss 0.017112f
C1764 avdd.n253 dvss 0.024064f
C1765 avdd.n254 dvss 0.022994f
C1766 avdd.n255 dvss 0.014552f
C1767 avdd.n256 dvss 0.017112f
C1768 avdd.t53 dvss 0.059823f
C1769 avdd.n261 dvss 0.012834f
C1770 avdd.n262 dvss 0.014552f
C1771 avdd.n263 dvss 0.077636f
C1772 avdd.n264 dvss 0.014552f
C1773 avdd.n265 dvss 0.017112f
C1774 avdd.n266 dvss 0.028342f
C1775 avdd.n269 dvss 0.062316f
C1776 avdd.n273 dvss 0.014552f
C1777 avdd.n274 dvss 0.015508f
C1778 avdd.n275 dvss 0.024598f
C1779 avdd.n278 dvss 0.034754f
C1780 avdd.n279 dvss 0.039051f
C1781 avdd.t35 dvss 0.01586f
C1782 avdd.n280 dvss 0.059429f
C1783 avdd.t50 dvss 0.01586f
C1784 avdd.n281 dvss 0.059429f
C1785 avdd.n282 dvss 0.017112f
C1786 avdd.n283 dvss 0.012834f
C1787 avdd.n286 dvss 0.16858f
C1788 avdd.t34 dvss 0.169991f
C1789 avdd.n287 dvss 0.077271f
C1790 avdd.t55 dvss 0.059823f
C1791 avdd.n288 dvss 0.097213f
C1792 avdd.t40 dvss 0.059823f
C1793 avdd.n289 dvss 0.079764f
C1794 avdd.n292 dvss 0.024064f
C1795 avdd.n293 dvss 0.014552f
C1796 avdd.n294 dvss 0.077636f
C1797 avdd.n295 dvss 0.012834f
C1798 avdd.n296 dvss 0.017112f
C1799 avdd.n297 dvss 0.077635f
C1800 avdd.n298 dvss 0.014438f
C1801 avdd.n299 dvss 0.018716f
C1802 avdd.n303 dvss 0.09472f
C1803 avdd.t42 dvss 0.059823f
C1804 avdd.n304 dvss 0.084749f
C1805 avdd.n305 dvss 0.097213f
C1806 avdd.t68 dvss 0.059823f
C1807 avdd.n306 dvss 0.072286f
C1808 avdd.n310 dvss 0.012834f
C1809 avdd.n311 dvss 0.017112f
C1810 avdd.n312 dvss 0.077635f
C1811 avdd.n313 dvss 0.017112f
C1812 avdd.n314 dvss 0.029946f
C1813 avdd.n315 dvss 0.017112f
C1814 avdd.n316 dvss 0.014552f
C1815 avdd.n317 dvss 0.077636f
C1816 avdd.n318 dvss 0.012834f
C1817 avdd.n319 dvss 0.014552f
C1818 avdd.n320 dvss 0.077635f
C1819 avdd.n321 dvss 0.017112f
C1820 avdd.n322 dvss 0.012834f
C1821 avdd.n325 dvss 0.069794f
C1822 avdd.n326 dvss 0.087242f
C1823 avdd.t44 dvss 0.059823f
C1824 avdd.n327 dvss 0.064808f
C1825 avdd.n328 dvss 0.092227f
C1826 avdd.n331 dvss 0.027272f
C1827 avdd.n332 dvss 0.019786f
C1828 avdd.n334 dvss 0.077635f
C1829 avdd.n335 dvss 0.017112f
C1830 avdd.n336 dvss 0.012834f
C1831 avdd.n339 dvss 0.097213f
C1832 avdd.t62 dvss 0.059823f
C1833 avdd.n340 dvss 0.077271f
C1834 avdd.n341 dvss 0.079764f
C1835 avdd.n344 dvss 0.097213f
C1836 avdd.t64 dvss 0.059823f
C1837 avdd.n345 dvss 0.062316f
C1838 avdd.n346 dvss 0.09472f
C1839 avdd.t32 dvss 0.059823f
C1840 avdd.n347 dvss 0.084749f
C1841 avdd.n349 dvss 0.072286f
C1842 avdd.t38 dvss 0.059823f
C1843 avdd.n350 dvss 0.097213f
C1844 avdd.t36 dvss 0.059823f
C1845 avdd.n351 dvss 0.069794f
C1846 avdd.n353 dvss 0.087242f
C1847 avdd.t51 dvss 0.059823f
C1848 avdd.n354 dvss 0.092227f
C1849 avdd.n355 dvss 0.064808f
C1850 avdd.t48 dvss 0.189627f
C1851 avdd.n356 dvss 0.071768f
C1852 avdd.n357 dvss 0.017112f
C1853 avdd.t58 dvss 0.015885f
C1854 avdd.n358 dvss 0.054551f
C1855 avdd.t49 dvss 0.015885f
C1856 avdd.n359 dvss 0.054551f
C1857 avdd.n361 dvss 0.012834f
C1858 avdd.n365 dvss 0.027272f
C1859 avdd.n366 dvss 0.017112f
C1860 avdd.n367 dvss 0.077635f
C1861 avdd.n368 dvss 0.017112f
C1862 avdd.n369 dvss 0.012834f
C1863 avdd.n372 dvss 0.029946f
C1864 avdd.n373 dvss 0.017112f
C1865 avdd.n374 dvss 0.077635f
C1866 avdd.n375 dvss 0.017112f
C1867 avdd.n376 dvss 0.012834f
C1868 avdd.n380 dvss 0.018181f
C1869 avdd.n381 dvss 1.62649f
C1870 avdd.n382 dvss 1.55534f
C1871 avdd.t25 dvss 16.3671f
C1872 avdd.t121 dvss 26.856901f
C1873 avdd.n383 dvss 4.72394f
C1874 avdd.n384 dvss 2.89188f
C1875 avdd.t99 dvss 4.24911f
C1876 avdd.t122 dvss 6.65055f
C1877 avdd.n385 dvss 2.73115f
C1878 avdd.t93 dvss 0.033086f
C1879 avdd.t29 dvss 0.031855f
C1880 avdd.n386 dvss 0.018062f
C1881 avdd.n387 dvss 0.306499f
C1882 avdd.n388 dvss 0.018068f
C1883 avdd.n389 dvss 0.155315f
C1884 avdd.n390 dvss 0.018056f
C1885 avdd.n391 dvss 0.154309f
C1886 avdd.t7 dvss 0.03146f
C1887 avdd.n392 dvss 0.138002f
C1888 avdd.n393 dvss 0.688157f
C1889 avdd.n394 dvss 0.079462f
C1890 avdd.n395 dvss 0.080116f
C1891 avdd.n396 dvss 0.357245f
C1892 avdd.n397 dvss 0.357405f
C1893 avdd.t113 dvss 0.139734f
C1894 avdd.n398 dvss 0.020098f
C1895 avdd.t97 dvss 0.311517f
C1896 avdd.n399 dvss 0.044621f
C1897 avdd.n400 dvss 0.035523f
C1898 avdd.n401 dvss 0.026448f
C1899 avdd.n402 dvss 0.021115f
C1900 avdd.n403 dvss 0.03085f
C1901 avdd.n404 dvss 0.046523f
C1902 avdd.n405 dvss 0.062878f
C1903 avdd.n406 dvss 0.041845f
C1904 avdd.n407 dvss 0.018666f
C1905 avdd.n408 dvss 0.011781f
C1906 avdd.n409 dvss 0.027563f
C1907 avdd.n410 dvss 0.037102f
C1908 avdd.n411 dvss 0.024876f
C1909 avdd.n412 dvss 0.02162f
C1910 avdd.t6 dvss 0.317932f
C1911 avdd.n413 dvss 0.279468f
C1912 avdd.t82 dvss 0.311517f
C1913 avdd.t4 dvss 0.311517f
C1914 avdd.n414 dvss 0.279468f
C1915 avdd.t86 dvss 0.311517f
C1916 avdd.t92 dvss 0.279468f
C1917 avdd.n415 dvss 0.036975f
C1918 avdd.n416 dvss 0.035523f
C1919 avdd.n417 dvss 0.020098f
C1920 avdd.n418 dvss 0.011781f
C1921 avdd.n419 dvss 0.038183f
C1922 avdd.n420 dvss 0.024876f
C1923 avdd.n421 dvss 0.064683f
C1924 avdd.n422 dvss 0.041845f
C1925 avdd.t28 dvss 0.326003f
C1926 avdd.n423 dvss 0.279468f
C1927 avdd.t84 dvss 0.311517f
C1928 avdd.t96 dvss 0.279468f
C1929 avdd.n424 dvss 0.036975f
C1930 avdd.n425 dvss 0.02162f
C1931 avdd.n426 dvss 0.021115f
C1932 avdd.n427 dvss 0.018666f
C1933 avdd.n428 dvss 0.03085f
C1934 avdd.n429 dvss 0.279468f
C1935 avdd.t100 dvss 0.282032f
C1936 avdd.n430 dvss 0.169219f
C1937 avdd.n431 dvss 0.115351f
C1938 avdd.n432 dvss 0.204694f
C1939 avdd.n433 dvss 0.357597f
C1940 avdd.n434 dvss 1.79539f
C1941 avdd.n435 dvss 1.26028f
C1942 avdd.n436 dvss 2.59575f
C1943 avdd.n437 dvss 4.36713f
C1944 avdd.n438 dvss 1.22699f
C1945 avdd.n439 dvss 1.82106f
C1946 avdd.n440 dvss 1.50595f
C1947 avdd.n441 dvss 1.52061f
C1948 avdd.n442 dvss 1.38908f
C1949 avdd.n443 dvss 1.32158f
C1950 avdd.n444 dvss 0.597165f
C1951 avdd.n445 dvss 1.01141f
C1952 avdd.n446 dvss 2.18305f
C1953 avdd.n447 dvss 0.890124f
C1954 avdd.n448 dvss 0.759271f
C1955 avdd.n449 dvss 3.94452f
C1956 avdd.n450 dvss 7.45013f
C1957 avdd.n451 dvss 6.12291f
C1958 avdd.n452 dvss 0.907843f
C1959 avdd.n453 dvss 1.83885f
C1960 avdd.n454 dvss 2.1652f
C1961 avdd.n455 dvss 1.92115f
C1962 avdd.n456 dvss 3.40097f
C1963 avdd.n457 dvss 1.66906f
C1964 avdd.n458 dvss 0.619763f
C1965 avdd.n459 dvss 1.0259f
C1966 avdd.n460 dvss 0.176937f
C1967 avdd.n461 dvss 0.349251f
C1968 avdd.n462 dvss 0.086572f
C1969 avdd.n463 dvss 0.014431f
C1970 avdd.n464 dvss 0.167396f
C1971 avdd.t117 dvss 0.014999f
C1972 avdd.n465 dvss 0.064301f
C1973 avdd.n466 dvss 0.058637f
C1974 avdd.n467 dvss 0.058637f
C1975 avdd.t116 dvss 0.637448f
C1976 avdd.t20 dvss 1.62336f
C1977 avdd.n468 dvss 0.07071f
C1978 avdd.n469 dvss 0.022579f
C1979 avdd.n470 dvss 0.04826f
C1980 avdd.n471 dvss 0.035296f
C1981 avdd.t110 dvss 0.014999f
C1982 avdd.n473 dvss 0.45767f
C1983 avdd.n474 dvss 0.078493f
C1984 avdd.n475 dvss 0.051564f
C1985 avdd.n476 dvss 0.04826f
C1986 avdd.n477 dvss 0.07071f
C1987 avdd.n478 dvss 0.033554f
C1988 avdd.n479 dvss 0.049998f
C1989 avdd.n480 dvss 0.602406f
C1990 avdd.n481 dvss 0.040477f
C1991 avdd.n482 dvss 0.057854f
C1992 avdd.n483 dvss 0.057854f
C1993 avdd.n484 dvss 0.058637f
C1994 avdd.n486 dvss 0.483436f
C1995 avdd.n487 dvss 0.150155f
C1996 avdd.n488 dvss 0.286525f
C1997 avdd.n489 dvss 0.379085f
C1998 avdd.n490 dvss 0.058637f
C1999 avdd.t118 dvss 0.653542f
C2000 avdd.n491 dvss 0.637448f
C2001 avdd.n492 dvss 0.022579f
C2002 avdd.t119 dvss 0.014999f
C2003 avdd.n493 dvss 0.03558f
C2004 avdd.n494 dvss 0.033251f
C2005 avdd.n495 dvss 0.026884f
C2006 avdd.n496 dvss 0.018588f
C2007 avdd.n498 dvss 0.071052f
C2008 avdd.n499 dvss 0.064914f
C2009 avdd.n500 dvss 0.026472f
C2010 avdd.n501 dvss 0.046564f
C2011 avdd.n502 dvss 0.04826f
C2012 avdd.n503 dvss 0.648557f
C2013 avdd.n504 dvss 0.047477f
C2014 avdd.n505 dvss 0.110862f
C2015 avdd.n506 dvss 0.198254f
C2016 avdd.n507 dvss 0.495986f
C2017 avdd.n508 dvss 0.196241f
C2018 avdd.n509 dvss 0.297794f
C2019 avdd.n510 dvss 0.087115f
C2020 avdd.n511 dvss 0.089258f
C2021 avdd.n512 dvss 0.08289f
C2022 avdd.n513 dvss 0.047477f
C2023 avdd.n514 dvss 0.648557f
C2024 avdd.n515 dvss 0.022579f
C2025 avdd.n516 dvss 0.038328f
C2026 avdd.n517 dvss 0.054238f
C2027 avdd.n518 dvss 0.026472f
C2028 avdd.n519 dvss 0.046564f
C2029 avdd.n520 dvss 0.04826f
C2030 avdd.n521 dvss 0.047477f
C2031 avdd.n522 dvss 0.477237f
C2032 avdd.n523 dvss 0.477237f
C2033 avdd.n524 dvss 0.072374f
C2034 avdd.n525 dvss 0.010973f
C2035 avdd.n526 dvss 0.016209f
C2036 avdd.n528 dvss 0.18742f
C2037 avdd.n529 dvss 0.087461f
C2038 avdd.n530 dvss 0.029454f
C2039 avdd.n531 dvss 0.339309f
C2040 avdd.n532 dvss 0.17581f
C2041 avdd.n533 dvss 0.253072f
C2042 avdd.n534 dvss 0.299937f
C2043 avdd.n535 dvss 1.33435f
C2044 avdd.n536 dvss 2.35062f
C2045 avdd.n537 dvss 0.834531f
C2046 porb_h[0].t2 dvss 0.015362f
C2047 porb_h[0].t15 dvss 0.015362f
C2048 porb_h[0].n0 dvss 0.063194f
C2049 porb_h[0].t21 dvss 0.030725f
C2050 porb_h[0].t20 dvss 0.030725f
C2051 porb_h[0].n1 dvss 0.07289f
C2052 porb_h[0].n2 dvss 0.233605f
C2053 porb_h[0].n3 dvss 0.018072f
C2054 porb_h[0].n4 dvss 0.016942f
C2055 porb_h[0].n5 dvss 0.125833f
C2056 porb_h[0].t9 dvss 0.015362f
C2057 porb_h[0].t8 dvss 0.015362f
C2058 porb_h[0].n6 dvss 0.063195f
C2059 porb_h[0].t30 dvss 0.030725f
C2060 porb_h[0].t29 dvss 0.030725f
C2061 porb_h[0].n7 dvss 0.07289f
C2062 porb_h[0].n8 dvss 0.233605f
C2063 porb_h[0].n9 dvss 0.205156f
C2064 porb_h[0].t4 dvss 0.015362f
C2065 porb_h[0].t14 dvss 0.015362f
C2066 porb_h[0].n10 dvss 0.063195f
C2067 porb_h[0].t26 dvss 0.030725f
C2068 porb_h[0].t25 dvss 0.030725f
C2069 porb_h[0].n11 dvss 0.07289f
C2070 porb_h[0].n12 dvss 0.233605f
C2071 porb_h[0].n13 dvss 0.229283f
C2072 porb_h[0].t5 dvss 0.015362f
C2073 porb_h[0].t13 dvss 0.015362f
C2074 porb_h[0].n14 dvss 0.063195f
C2075 porb_h[0].t28 dvss 0.030725f
C2076 porb_h[0].t24 dvss 0.030725f
C2077 porb_h[0].n15 dvss 0.07289f
C2078 porb_h[0].n16 dvss 0.233605f
C2079 porb_h[0].n17 dvss 0.229283f
C2080 porb_h[0].t0 dvss 0.015362f
C2081 porb_h[0].t6 dvss 0.015362f
C2082 porb_h[0].n18 dvss 0.063195f
C2083 porb_h[0].t19 dvss 0.030725f
C2084 porb_h[0].t27 dvss 0.030725f
C2085 porb_h[0].n19 dvss 0.07289f
C2086 porb_h[0].n20 dvss 0.233605f
C2087 porb_h[0].n21 dvss 0.229283f
C2088 porb_h[0].t7 dvss 0.015362f
C2089 porb_h[0].t1 dvss 0.015362f
C2090 porb_h[0].n22 dvss 0.063195f
C2091 porb_h[0].t22 dvss 0.030725f
C2092 porb_h[0].t17 dvss 0.030725f
C2093 porb_h[0].n23 dvss 0.07289f
C2094 porb_h[0].n24 dvss 0.233605f
C2095 porb_h[0].n25 dvss 0.229283f
C2096 porb_h[0].t3 dvss 0.015362f
C2097 porb_h[0].t11 dvss 0.015362f
C2098 porb_h[0].n26 dvss 0.063195f
C2099 porb_h[0].t18 dvss 0.030725f
C2100 porb_h[0].t23 dvss 0.030725f
C2101 porb_h[0].n27 dvss 0.07289f
C2102 porb_h[0].n28 dvss 0.233605f
C2103 porb_h[0].n29 dvss 0.229283f
C2104 porb_h[0].t12 dvss 0.015362f
C2105 porb_h[0].t10 dvss 0.015362f
C2106 porb_h[0].n30 dvss 0.063195f
C2107 porb_h[0].t16 dvss 0.030725f
C2108 porb_h[0].t31 dvss 0.030725f
C2109 porb_h[0].n31 dvss 0.07289f
C2110 porb_h[0].n32 dvss 0.233605f
C2111 porb_h[0].n33 dvss 0.433858f
C2112 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n0 dvss 2.54524f
C2113 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n1 dvss 1.79517f
C2114 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n2 dvss 0.090207f
C2115 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n3 dvss 0.10921f
C2116 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n4 dvss 0.018812f
C2117 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n5 dvss 0.119127f
C2118 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n6 dvss 0.119093f
C2119 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n7 dvss 0.018812f
C2120 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n8 dvss 0.119127f
C2121 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n9 dvss 0.119093f
C2122 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n10 dvss 0.119127f
C2123 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n11 dvss 0.119093f
C2124 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n12 dvss 0.018812f
C2125 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n13 dvss 0.119127f
C2126 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n14 dvss 0.119093f
C2127 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n15 dvss 0.119127f
C2128 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n16 dvss 0.119093f
C2129 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n17 dvss 0.119127f
C2130 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n18 dvss 0.100089f
C2131 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n19 dvss 0.10921f
C2132 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n20 dvss 0.119127f
C2133 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n21 dvss 0.119093f
C2134 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n22 dvss 0.018812f
C2135 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n23 dvss 0.119127f
C2136 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n24 dvss 0.119093f
C2137 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n25 dvss 0.119127f
C2138 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n26 dvss 0.119093f
C2139 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n27 dvss 0.018812f
C2140 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n28 dvss 0.119127f
C2141 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n29 dvss 0.119093f
C2142 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n30 dvss 0.119127f
C2143 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n31 dvss 0.119093f
C2144 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n32 dvss 0.119127f
C2145 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n33 dvss 0.100089f
C2146 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n34 dvss 0.090207f
C2147 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n35 dvss 2.12882f
C2148 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n36 dvss 0.018812f
C2149 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n37 dvss 0.018812f
C2150 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n38 dvss 0.018812f
C2151 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n39 dvss 0.018812f
C2152 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n40 dvss 0.018812f
C2153 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n41 dvss 0.018812f
C2154 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n42 dvss 0.018812f
C2155 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t21 dvss 0.043796f
C2156 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t55 dvss 0.098823f
C2157 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t18 dvss 0.053679f
C2158 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t46 dvss 0.10355f
C2159 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n43 dvss 0.110577f
C2160 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t30 dvss 0.098823f
C2161 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t51 dvss 0.043796f
C2162 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t54 dvss 0.098823f
C2163 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t20 dvss 0.043796f
C2164 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t63 dvss 0.043796f
C2165 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t31 dvss 0.098823f
C2166 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t27 dvss 0.043796f
C2167 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t4 dvss 0.098823f
C2168 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t38 dvss 0.098823f
C2169 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t67 dvss 0.043796f
C2170 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t14 dvss 0.098823f
C2171 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t35 dvss 0.043796f
C2172 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t13 dvss 0.043796f
C2173 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t49 dvss 0.098823f
C2174 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t37 dvss 0.043796f
C2175 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t16 dvss 0.098823f
C2176 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t15 dvss 0.098823f
C2177 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t43 dvss 0.043796f
C2178 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t48 dvss 0.098823f
C2179 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t12 dvss 0.043796f
C2180 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t24 dvss 0.043796f
C2181 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t58 dvss 0.098823f
C2182 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t23 dvss 0.043796f
C2183 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t57 dvss 0.098823f
C2184 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n44 dvss 0.026757f
C2185 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t32 dvss 0.098823f
C2186 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t56 dvss 0.043796f
C2187 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t6 dvss 0.053642f
C2188 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t33 dvss 0.108644f
C2189 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n45 dvss 0.10592f
C2190 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n46 dvss 0.026861f
C2191 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n47 dvss 0.026899f
C2192 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n48 dvss 0.025223f
C2193 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t0 dvss 0.049857f
C2194 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t1 dvss 0.04919f
C2195 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t3 dvss 0.032567f
C2196 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t2 dvss 0.032567f
C2197 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n49 dvss 0.06859f
C2198 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t62 dvss 0.043796f
C2199 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t8 dvss 0.098823f
C2200 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t60 dvss 0.10355f
C2201 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t59 dvss 0.053679f
C2202 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n50 dvss 0.110581f
C2203 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t39 dvss 0.098823f
C2204 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t34 dvss 0.043796f
C2205 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t7 dvss 0.098823f
C2206 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t61 dvss 0.043796f
C2207 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t40 dvss 0.043796f
C2208 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t41 dvss 0.098823f
C2209 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t9 dvss 0.043796f
C2210 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t17 dvss 0.098823f
C2211 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t50 dvss 0.098823f
C2212 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t42 dvss 0.043796f
C2213 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t25 dvss 0.098823f
C2214 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t19 dvss 0.043796f
C2215 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t53 dvss 0.043796f
C2216 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t65 dvss 0.098823f
C2217 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t22 dvss 0.043796f
C2218 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t29 dvss 0.098823f
C2219 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t28 dvss 0.098823f
C2220 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t26 dvss 0.043796f
C2221 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t64 dvss 0.098823f
C2222 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t52 dvss 0.043796f
C2223 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t5 dvss 0.043796f
C2224 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t11 dvss 0.098823f
C2225 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t66 dvss 0.043796f
C2226 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t10 dvss 0.098823f
C2227 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n51 dvss 0.026757f
C2228 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t44 dvss 0.098823f
C2229 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t36 dvss 0.043796f
C2230 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t47 dvss 0.108644f
C2231 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.t45 dvss 0.053642f
C2232 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n52 dvss 0.10592f
C2233 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n53 dvss 0.026861f
C2234 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n54 dvss 0.026899f
C2235 x2.por_output_driver_h_0/sky130_fd_sc_hvl__inv_16_0.A.n55 dvss 0.025223f
C2236 avss.n1 dvss 0.037248f
C2237 avss.n2 dvss 0.028216f
C2238 avss.n4 dvss 0.011049f
C2239 avss.n9 dvss 0.029585f
C2240 avss.n10 dvss 0.037559f
C2241 avss.n11 dvss 0.015761f
C2242 avss.n19 dvss 0.089809f
C2243 avss.n20 dvss 0.029376f
C2244 avss.n24 dvss 0.033971f
C2245 avss.t72 dvss 0.050394f
C2246 avss.n28 dvss 0.018361f
C2247 avss.n29 dvss 0.131469f
C2248 avss.n30 dvss 0.07762f
C2249 avss.n32 dvss 0.015102f
C2250 avss.t20 dvss 0.125958f
C2251 avss.t31 dvss 0.046435f
C2252 avss.n35 dvss 0.012328f
C2253 avss.n39 dvss 0.045302f
C2254 avss.n40 dvss 0.048151f
C2255 avss.t24 dvss 0.031721f
C2256 avss.n41 dvss 0.012682f
C2257 avss.t25 dvss 0.046919f
C2258 avss.n44 dvss 0.012748f
C2259 avss.n46 dvss 0.011651f
C2260 avss.n49 dvss 0.012619f
C2261 avss.n55 dvss 0.025996f
C2262 avss.t3 dvss 0.043141f
C2263 avss.n58 dvss 0.015658f
C2264 avss.n59 dvss 0.015638f
C2265 avss.n63 dvss 0.046671f
C2266 avss.n65 dvss 0.022108f
C2267 avss.n72 dvss 0.032252f
C2268 avss.n73 dvss 0.045289f
C2269 avss.n74 dvss 0.028282f
C2270 avss.n77 dvss 0.038792f
C2271 avss.t59 dvss 0.035925f
C2272 avss.n79 dvss 0.014041f
C2273 avss.t53 dvss 0.020016f
C2274 avss.t45 dvss 0.046435f
C2275 avss.t33 dvss 0.029428f
C2276 avss.n85 dvss 0.031721f
C2277 avss.t27 dvss 0.046435f
C2278 avss.n93 dvss 0.029683f
C2279 avss.n94 dvss 0.034768f
C2280 avss.n100 dvss 0.039107f
C2281 avss.n101 dvss 0.034802f
C2282 avss.n111 dvss 0.03254f
C2283 avss.n116 dvss 0.02415f
C2284 avss.n117 dvss 0.026557f
C2285 avss.n118 dvss 0.032102f
C2286 avss.t66 dvss 0.033802f
C2287 avss.n135 dvss 0.062375f
C2288 avss.n136 dvss 0.213542f
C2289 avss.t15 dvss 0.076802f
C2290 avss.n140 dvss 0.0118f
C2291 avss.t46 dvss 0.046197f
C2292 avss.n141 dvss 0.028733f
C2293 avss.n142 dvss 0.029162f
C2294 avss.t44 dvss 0.048744f
C2295 avss.t47 dvss 0.04874f
C2296 avss.t12 dvss 0.04874f
C2297 avss.t30 dvss 0.04874f
C2298 avss.t61 dvss 0.04874f
C2299 avss.t74 dvss 0.04874f
C2300 avss.n145 dvss 0.031721f
C2301 avss.t60 dvss 0.032868f
C2302 avss.t68 dvss 0.064039f
C2303 avss.t71 dvss 0.049384f
C2304 avss.t28 dvss 0.04874f
C2305 avss.t41 dvss 0.04874f
C2306 avss.n149 dvss 0.060317f
C2307 avss.n150 dvss 0.073481f
C2308 avss.n152 dvss 0.012971f
C2309 avss.n154 dvss 0.015617f
C2310 avss.n158 dvss 0.116928f
C2311 avss.n159 dvss 0.060543f
C2312 avss.n160 dvss 0.502919f
C2313 avss.n161 dvss 0.011551f
C2314 avss.n162 dvss 0.011551f
C2315 avss.n163 dvss 0.035703f
C2316 avss.n165 dvss 0.029383f
C2317 avss.n166 dvss 0.832393f
C2318 avss.n167 dvss 0.293502f
C2319 avss.n168 dvss 0.018865f
C2320 avss.n169 dvss 0.01305f
C2321 avss.n170 dvss 0.011551f
C2322 avss.n171 dvss 0.039985f
C2323 avss.n172 dvss 0.011523f
C2324 avss.n173 dvss 0.512701f
C2325 avss.n174 dvss 0.011551f
C2326 avss.n175 dvss 0.234778f
C2327 avss.n176 dvss 0.043567f
C2328 avss.n180 dvss 0.148592f
C2329 avss.n185 dvss 0.011542f
C2330 avss.n190 dvss 0.019234f
C2331 avss.n191 dvss 0.019234f
C2332 avss.n200 dvss 0.014308f
C2333 avss.n211 dvss 0.013099f
C2334 avss.n212 dvss 0.013928f
C2335 avss.n213 dvss 0.023186f
C2336 avss.n214 dvss 0.010412f
C2337 avss.n215 dvss 0.066217f
C2338 avss.n216 dvss 0.040949f
C2339 avss.n217 dvss 0.142861f
C2340 avss.n218 dvss 0.291589f
C2341 avss.n219 dvss 0.06632f
C2342 avss.n220 dvss 0.245902f
C2343 avss.n222 dvss 0.021541f
C2344 avss.n230 dvss 0.074589f
C2345 avss.n231 dvss 0.068598f
C2346 avss.n232 dvss 0.159539f
C2347 avss.n238 dvss 0.03272f
C2348 avss.n342 dvss 0.063367f
C2349 avss.n397 dvss 0.049001f
C2350 avss.n398 dvss 0.081511f
C2351 avss.n477 dvss 0.08045f
C2352 avss.n499 dvss 0.023308f
C2353 avss.n500 dvss 0.061411f
C2354 avss.n505 dvss 0.116349f
C2355 avss.n506 dvss 0.173033f
C2356 avss.n511 dvss 0.03482f
C2357 avss.n516 dvss 0.01518f
C2358 avss.n517 dvss 0.031996f
C2359 avss.n525 dvss 0.01741f
C2360 avss.n533 dvss 0.022218f
C2361 avss.n534 dvss 0.03482f
C2362 avss.n541 dvss 0.062841f
C2363 avss.n542 dvss 0.102379f
C2364 avss.n543 dvss 0.127921f
C2365 avss.n546 dvss 0.050336f
C2366 avss.n551 dvss 0.154605f
C2367 avss.n552 dvss 0.066947f
C2368 avss.n553 dvss 0.059893f
C2369 avss.n555 dvss 0.048584f
C2370 avss.n565 dvss 0.048584f
C2371 avss.n580 dvss 0.048584f
C2372 avss.n581 dvss 0.038047f
C2373 avss.n582 dvss 0.024292f
C2374 avss.n583 dvss 0.034668f
C2375 avss.n587 dvss 0.019862f
C2376 avss.n588 dvss 0.01508f
C2377 avss.n593 dvss 0.026786f
C2378 avss.n594 dvss 0.023246f
C2379 avss.n597 dvss 0.04642f
C2380 avss.n601 dvss 0.045418f
C2381 avss.n602 dvss 0.057041f
C2382 avss.n615 dvss 0.027238f
C2383 avss.n620 dvss 0.019758f
C2384 avss.n622 dvss 0.024403f
C2385 avss.n623 dvss 0.016547f
C2386 avss.n627 dvss 0.023422f
C2387 avss.n631 dvss 0.010502f
C2388 avss.n632 dvss 0.036206f
C2389 avss.n633 dvss 0.057869f
C2390 avss.n653 dvss 0.02762f
C2391 avss.n658 dvss 0.439971f
C2392 avss.n659 dvss 0.045005f
C2393 avss.n732 dvss 0.036224f
C2394 avss.n733 dvss 0.032084f
C2395 avss.n741 dvss 0.028112f
C2396 avss.n745 dvss 0.024139f
C2397 avss.n753 dvss 0.024139f
C2398 avss.n754 dvss 0.029792f
C2399 avss.n761 dvss 0.02618f
C2400 avss.n768 dvss 0.064819f
C2401 avss.n782 dvss 0.035445f
C2402 avss.n783 dvss 0.035445f
C2403 avss.n789 dvss 0.024139f
C2404 avss.n797 dvss 0.024139f
C2405 avss.n798 dvss 0.024139f
C2406 avss.n805 dvss 0.08535f
C2407 avss.n806 dvss 0.081928f
C2408 avss.n809 dvss 0.028575f
C2409 avss.n810 dvss 0.022275f
C2410 avss.n811 dvss 0.110822f
C2411 avss.n812 dvss 0.104099f
C2412 avss.n814 dvss 0.033938f
C2413 avss.n815 dvss 0.032498f
C2414 avss.n819 dvss 0.017003f
C2415 avss.n874 dvss 0.016888f
C2416 avss.n875 dvss 0.068219f
C2417 avss.n876 dvss 0.041416f
C2418 avss.n877 dvss 0.019788f
C2419 avss.n889 dvss 0.068026f
C2420 avss.n890 dvss 0.290549f
C2421 avss.n891 dvss 0.117231f
C2422 avss.n892 dvss 0.129832f
C2423 avss.n893 dvss 0.049135f
C2424 avss.n894 dvss 0.094423f
C2425 avss.n901 dvss 0.068167f
C2426 avss.n911 dvss 0.095251f
C2427 avss.n912 dvss 0.04191f
C2428 avss.n919 dvss 0.08175f
C2429 avss.n920 dvss 0.079749f
C2430 avss.n921 dvss 0.035036f
C2431 avss.n922 dvss 0.019339f
C2432 avss.n936 dvss 0.013099f
C2433 avss.n940 dvss 0.031021f
C2434 avss.n941 dvss 1.30497f
C2435 avss.n942 dvss 0.789343f
C2436 avss.n943 dvss 1.0423f
C2437 avss.n944 dvss 0.789343f
C2438 avss.n945 dvss 0.784291f
C2439 avss.n946 dvss 0.789343f
C2440 avss.n947 dvss 0.784291f
C2441 avss.n948 dvss 0.789343f
C2442 avss.n949 dvss 0.784291f
C2443 avss.n950 dvss 0.789343f
C2444 avss.n951 dvss 0.784291f
C2445 avss.n952 dvss 0.789343f
C2446 avss.n953 dvss 0.784291f
C2447 avss.n954 dvss 0.789343f
C2448 avss.n955 dvss 0.784291f
C2449 avss.n956 dvss 0.789343f
C2450 avss.n957 dvss 0.784291f
C2451 avss.n958 dvss 0.789343f
C2452 avss.n959 dvss 0.739289f
C2453 avss.n960 dvss 1.30497f
C2454 avss.n961 dvss 0.789343f
C2455 avss.n962 dvss 1.0423f
C2456 avss.n963 dvss 0.789343f
C2457 avss.n964 dvss 0.784291f
C2458 avss.n965 dvss 0.789343f
C2459 avss.n966 dvss 0.784291f
C2460 avss.n967 dvss 0.789343f
C2461 avss.n968 dvss 0.784291f
C2462 avss.n969 dvss 0.789343f
C2463 avss.n970 dvss 0.784291f
C2464 avss.n971 dvss 0.789343f
C2465 avss.n972 dvss 0.784291f
C2466 avss.n973 dvss 0.789343f
C2467 avss.n974 dvss 0.784291f
C2468 avss.n975 dvss 0.789343f
C2469 avss.n976 dvss 0.784291f
C2470 avss.n977 dvss 0.789343f
C2471 avss.n978 dvss -3.27748f
C2472 avss.n979 dvss 1.30497f
C2473 avss.n980 dvss 0.789343f
C2474 avss.n981 dvss 1.0423f
C2475 avss.n982 dvss 0.789343f
C2476 avss.n983 dvss 0.784291f
C2477 avss.n984 dvss 0.789343f
C2478 avss.n985 dvss 0.784291f
C2479 avss.n986 dvss 0.789343f
C2480 avss.n987 dvss 0.784291f
C2481 avss.n988 dvss 0.789343f
C2482 avss.n989 dvss 0.784291f
C2483 avss.n990 dvss 0.789343f
C2484 avss.n991 dvss 0.784291f
C2485 avss.n992 dvss 0.789343f
C2486 avss.n993 dvss 0.784291f
C2487 avss.n994 dvss 0.789343f
C2488 avss.n995 dvss 0.784291f
C2489 avss.n996 dvss 0.789343f
C2490 avss.n997 dvss 0.750275f
C2491 avss.n998 dvss -13.5832f
C2492 avss.n999 dvss -8.493879f
C2493 avss.n1000 dvss 1.30497f
C2494 avss.n1001 dvss 0.789343f
C2495 avss.n1002 dvss 1.0423f
C2496 avss.n1003 dvss 0.789343f
C2497 avss.n1004 dvss 0.784291f
C2498 avss.n1005 dvss 0.789343f
C2499 avss.n1006 dvss 0.784291f
C2500 avss.n1007 dvss 0.789343f
C2501 avss.n1008 dvss 0.784291f
C2502 avss.n1009 dvss 0.789343f
C2503 avss.n1010 dvss 0.784291f
C2504 avss.n1011 dvss 0.789343f
C2505 avss.n1012 dvss 0.784291f
C2506 avss.n1013 dvss 0.789343f
C2507 avss.n1014 dvss 0.784291f
C2508 avss.n1015 dvss 0.789343f
C2509 avss.n1016 dvss 0.784291f
C2510 avss.n1017 dvss 0.789343f
C2511 avss.n1018 dvss -3.37571f
C2512 avss.n1019 dvss -4.29067f
C2513 avss.n1020 dvss 0.931146f
C2514 avss.n1021 dvss 0.396858f
C2515 avss.n1022 dvss 0.143298f
C2516 avss.n1023 dvss 0.180239f
C2517 avss.n1024 dvss 0.129016f
C2518 avss.n1025 dvss 0.227692f
C2519 avss.n1026 dvss 0.042252f
C2520 avss.n1027 dvss 0.049994f
C2521 avss.n1028 dvss 2.79876f
C2522 avss.n1029 dvss 4.72434f
C2523 avss.n1030 dvss 0.025697f
C2524 avss.n1031 dvss 0.089325f
C2525 avss.n1032 dvss 0.049729f
C2526 avss.n1033 dvss 3.3937f
C2527 avss.n1034 dvss 0.02041f
C2528 avss.n1035 dvss 0.062097f
C2529 avss.n1036 dvss 0.037279f
C2530 avss.n1037 dvss 0.036361f
C2531 avss.n1038 dvss 0.089861f
C2532 avss.n1039 dvss 0.114671f
C2533 avss.n1040 dvss 0.181236f
C2534 avss.n1041 dvss 0.088323f
C2535 avss.n1042 dvss 0.108534f
C2536 avss.n1043 dvss 0.03979f
C2537 avss.n1044 dvss 10.191401f
C2538 avss.n1045 dvss 4.69219f
C2539 avss.n1046 dvss 17.2493f
C2540 avss.n1047 dvss 0.057598f
C2541 avss.n1048 dvss 0.142503f
C2542 avss.n1049 dvss 0.150768f
C2543 avss.n1050 dvss 0.109138f
C2544 avss.n1051 dvss 0.114371f
C2545 avss.n1052 dvss 0.121994f
C2546 avss.n1053 dvss 0.105362f
C2547 avss.n1054 dvss 0.444556f
C2548 avss.n1055 dvss 0.46878f
C2549 avss.n1056 dvss -0.247953f
C2550 avss.n1057 dvss 0.061022f
C2551 avss.n1058 dvss 0.110534f
C2552 avss.n1059 dvss 0.016756f
C2553 avss.n1060 dvss 0.013222f
C2554 avss.n1063 dvss 0.085892f
C2555 avss.n1064 dvss 0.033379f
C2556 avss.n1070 dvss 0.084222f
C2557 avss.n1071 dvss 0.315383f
C2558 avss.n1072 dvss 0.38438f
C2559 avss.n1073 dvss 0.355553f
C2560 avss.n1074 dvss 0.010383f
C2561 avss.n1075 dvss 0.027814f
C2562 avss.n1076 dvss 0.087318f
C2563 avss.n1077 dvss 0.145205f
C2564 avss.n1078 dvss 0.013731f
C2565 avss.n1079 dvss 0.019413f
C2566 avss.n1080 dvss 0.407428f
C2567 avss.n1082 dvss 0.531422f
C2568 avss.n1084 dvss 0.012975f
C2569 avss.n1085 dvss 0.035695f
C2570 avss.n1086 dvss 0.011523f
C2571 avss.n1087 dvss 0.476832f
C2572 avss.n1088 dvss 0.632476f
C2573 avss.n1089 dvss 0.107466f
C2574 avss.n1090 dvss 0.098932f
C2575 avss.n1091 dvss 0.033219f
C2576 avss.n1095 dvss 0.020055f
C2577 avss.n1096 dvss 0.026371f
C2578 avss.n1100 dvss 0.020336f
C2579 avss.n1103 dvss 0.02733f
C2580 avss.n1104 dvss 0.017316f
C2581 avss.n1110 dvss 0.011674f
C2582 avss.t63 dvss 0.017875f
C2583 avss.n1115 dvss 0.011869f
C2584 avss.t9 dvss 0.039471f
C2585 avss.t1 dvss 0.039471f
C2586 avss.n1124 dvss 0.012275f
C2587 avss.n1131 dvss 0.010072f
C2588 avss.n1133 dvss 0.010557f
C2589 avss.t52 dvss 0.034979f
C2590 avss.n1145 dvss 0.016325f
C2591 avss.n1146 dvss 0.013855f
C2592 avss.n1147 dvss 0.013947f
C2593 avss.t65 dvss 0.053121f
C2594 avss.n1157 dvss 0.021119f
C2595 avss.n1158 dvss 0.01422f
C2596 avss.n1160 dvss 0.046435f
C2597 avss.t19 dvss 0.108148f
C2598 avss.n1167 dvss 0.036549f
C2599 avss.n1169 dvss 0.020292f
C2600 avss.n1175 dvss 0.018479f
C2601 avss.n1176 dvss 0.018479f
C2602 avss.t49 dvss 0.018479f
C2603 avss.n1192 dvss 0.033963f
C2604 avss.t18 dvss 0.018479f
C2605 avss.t48 dvss 0.018479f
C2606 avss.n1203 dvss 0.021695f
C2607 avss.n1204 dvss 0.027043f
C2608 avss.n1205 dvss 0.0175f
C2609 avss.n1206 dvss 0.013074f
C2610 avss.n1212 dvss 0.038357f
C2611 avss.n1213 dvss 0.028389f
C2612 avss.t17 dvss 0.031721f
C2613 avss.t58 dvss 0.053283f
C2614 avss.t39 dvss 0.053283f
C2615 avss.t70 dvss 0.058559f
C2616 avss.t56 dvss 0.062206f
C2617 avss.t23 dvss 0.04204f
C2618 avss.t0 dvss 0.059742f
C2619 avss.n1215 dvss 0.02525f
C2620 avss.n1217 dvss 0.033173f
C2621 avss.t7 dvss 0.041945f
C2622 avss.n1218 dvss 0.028708f
C2623 avss.n1223 dvss 0.012779f
C2624 avss.n1224 dvss 0.017401f
C2625 avss.n1225 dvss 0.013224f
C2626 avss.n1229 dvss 0.021402f
C2627 avss.t57 dvss 0.015861f
C2628 avss.t35 dvss 0.05246f
C2629 avss.t13 dvss 0.061925f
C2630 avss.t21 dvss 0.053124f
C2631 avss.t55 dvss 0.063443f
C2632 avss.t51 dvss 0.063443f
C2633 avss.t34 dvss 0.063443f
C2634 avss.t22 dvss 0.063443f
C2635 avss.t54 dvss 0.063443f
C2636 avss.t42 dvss 0.063443f
C2637 avss.t26 dvss 0.063443f
C2638 avss.t40 dvss 0.063443f
C2639 avss.t62 dvss 0.063443f
C2640 avss.t43 dvss 0.032486f
C2641 avss.n1231 dvss 0.038234f
C2642 avss.t38 dvss 0.062678f
C2643 avss.t75 dvss 0.051213f
C2644 avss.n1232 dvss 0.031721f
C2645 avss.t29 dvss 0.043951f
C2646 avss.t16 dvss 0.034206f
C2647 avss.n1233 dvss 0.025004f
C2648 avss.n1234 dvss 0.013842f
C2649 avss.t69 dvss 0.12005f
C2650 avss.n1241 dvss 0.028282f
C2651 avss.n1242 dvss 0.046435f
C2652 avss.n1244 dvss 0.014912f
C2653 avss.n1245 dvss 0.022984f
C2654 avss.n1246 dvss 0.040743f
C2655 avss.n1247 dvss 0.016268f
C2656 avss.n1248 dvss 0.067688f
C2657 avss.n1249 dvss 0.052779f
C2658 avss.n1250 dvss 0.033984f
C2659 avss.n1251 dvss 0.130675f
C2660 avss.n1252 dvss 0.027466f
C2661 avss.n1253 dvss 0.017246f
C2662 avss.n1255 dvss 1.15929f
C2663 avss.n1256 dvss 0.235246f
C2664 avss.t5 dvss 0.027591f
C2665 avss.n1260 dvss 0.013224f
C2666 avss.t32 dvss 0.034768f
C2667 avss.n1265 dvss 0.06528f
C2668 avss.n1266 dvss 0.068237f
C2669 avss.n1269 dvss 0.407873f
C2670 avss.n1270 dvss 0.348748f
C2671 a_5972_n290308.n0 dvss 1.90875f
C2672 a_5972_n290308.t5 dvss 1.10214f
C2673 a_5972_n290308.t4 dvss 0.048368f
C2674 a_5972_n290308.t0 dvss 0.096352f
C2675 a_5972_n290308.t1 dvss 0.09029f
C2676 a_5972_n290308.t3 dvss 1.10336f
C2677 a_5972_n290308.n1 dvss 1.62858f
C2678 a_5972_n290308.t2 dvss 0.222171f
C2679 x1.vbn.n0 dvss 1.32541f
C2680 x1.vbn.n1 dvss 0.711391f
C2681 x1.vbn.t5 dvss 0.413212f
C2682 x1.vbn.t4 dvss 0.405095f
C2683 x1.vbn.n2 dvss 0.698301f
C2684 x1.vbn.t8 dvss 0.405082f
C2685 x1.vbn.t10 dvss 0.413261f
C2686 x1.vbn.n3 dvss 0.648014f
C2687 x1.vbn.n4 dvss 0.512488f
C2688 x1.vbn.t6 dvss 0.175014f
C2689 x1.vbn.t3 dvss 0.222317f
C2690 x1.vbn.n5 dvss 1.21542f
C2691 x1.vbn.t1 dvss 0.407193f
C2692 x1.vbn.t0 dvss 0.054827f
C2693 x1.vbn.t2 dvss 0.093658f
C2694 x1.vbn.t7 dvss 0.4138f
C2695 x1.vbn.t9 dvss 0.405083f
C2696 x1.vbn.n6 dvss 0.629348f
C2697 a_4566_n291516.t3 dvss 0.336034f
C2698 a_4566_n291516.t2 dvss 0.050475f
C2699 a_4566_n291516.t1 dvss 1.22045f
C2700 a_4566_n291516.n0 dvss 0.916763f
C2701 a_4566_n291516.n1 dvss 1.56301f
C2702 a_4566_n291516.t0 dvss 0.213264f
C2703 x2.Td_L.n0 dvss 0.093879f
C2704 x2.Td_L.n1 dvss 0.559627f
C2705 x2.Td_L.n2 dvss 1.92623f
C2706 x2.Td_L.n3 dvss 0.116237f
C2707 x2.Td_L.n4 dvss 0.636203f
C2708 x2.Td_L.n5 dvss 0.119977f
C2709 x2.Td_L.t6 dvss 0.049756f
C2710 x2.Td_L.t12 dvss 0.049793f
C2711 x2.Td_L.n6 dvss 0.117398f
C2712 x2.Td_L.t7 dvss 0.045979f
C2713 x2.Td_L.t11 dvss 0.073839f
C2714 x2.Td_L.t10 dvss 0.127545f
C2715 x2.Td_L.t14 dvss 0.094244f
C2716 x2.Td_L.n7 dvss 0.117087f
C2717 x2.Td_L.n8 dvss 1.73539f
C2718 x2.Td_L.t13 dvss 0.049761f
C2719 x2.Td_L.n9 dvss 0.117404f
C2720 x2.Td_L.t8 dvss 0.049779f
C2721 x2.Td_L.n10 dvss 0.113872f
C2722 x2.Td_L.t9 dvss 0.047826f
C2723 x2.Td_L.t15 dvss 0.047866f
C2724 x2.Td_L.n11 dvss 0.1117f
C2725 x2.Td_L.t1 dvss 0.016025f
C2726 x2.Td_L.t0 dvss 0.016025f
C2727 x2.Td_L.n12 dvss 0.035099f
C2728 x2.Td_L.t2 dvss 0.022435f
C2729 x2.Td_L.t4 dvss 0.022435f
C2730 x2.Td_L.n13 dvss 0.047226f
C2731 x2.Td_L.t3 dvss 0.022435f
C2732 x2.Td_L.t5 dvss 0.022435f
C2733 x2.Td_L.n14 dvss 0.046487f
C2734 x2.Td_L.n15 dvss 0.532351f
C2735 a_32918_n290853.n0 dvss 0.410268f
C2736 a_32918_n290853.n1 dvss 0.543744f
C2737 a_32918_n290853.n2 dvss 0.679078f
C2738 a_32918_n290853.t1 dvss 0.047481f
C2739 a_32918_n290853.t0 dvss 0.034067f
C2740 a_32918_n290853.n3 dvss 0.077122f
C2741 a_32918_n290853.t5 dvss 0.031982f
C2742 a_32918_n290853.t8 dvss 0.032006f
C2743 a_32918_n290853.n4 dvss 0.075509f
C2744 a_32918_n290853.t3 dvss 0.031982f
C2745 a_32918_n290853.n5 dvss 0.075523f
C2746 a_32918_n290853.t6 dvss 0.032006f
C2747 a_32918_n290853.n6 dvss 0.075527f
C2748 a_32918_n290853.n7 dvss 0.073272f
C2749 a_32918_n290853.t7 dvss 0.030742f
C2750 a_32918_n290853.t4 dvss 0.030768f
C2751 a_32918_n290853.n8 dvss 0.071851f
C2752 a_32918_n290853.t2 dvss 0.047073f
C2753 a_37002_n287783.n0 dvss 0.686222f
C2754 a_37002_n287783.n1 dvss 1.02628f
C2755 a_37002_n287783.t3 dvss 0.022918f
C2756 a_37002_n287783.t1 dvss 0.033532f
C2757 a_37002_n287783.t0 dvss 0.033919f
C2758 a_37002_n287783.t5 dvss 0.163037f
C2759 a_37002_n287783.t4 dvss 0.09889f
C2760 a_37002_n287783.t7 dvss 0.16472f
C2761 a_37002_n287783.t6 dvss 0.09891f
C2762 a_37002_n287783.n2 dvss 0.048656f
C2763 a_37002_n287783.t2 dvss 0.022918f
C2764 a_36398_n287783.n0 dvss 0.647187f
C2765 a_36398_n287783.n1 dvss 1.26319f
C2766 a_36398_n287783.t2 dvss 0.023037f
C2767 a_36398_n287783.t7 dvss 0.163788f
C2768 a_36398_n287783.t5 dvss 0.09923f
C2769 a_36398_n287783.t6 dvss 0.163788f
C2770 a_36398_n287783.t4 dvss 0.09923f
C2771 a_36398_n287783.t3 dvss 0.033735f
C2772 a_36398_n287783.t1 dvss 0.034222f
C2773 a_36398_n287783.n2 dvss 0.049554f
C2774 a_36398_n287783.t0 dvss 0.023037f
C2775 a_25883_n288267.n0 dvss 0.041155f
C2776 a_25883_n288267.n1 dvss 0.02644f
C2777 a_25883_n288267.n2 dvss 0.26314f
C2778 a_25883_n288267.t0 dvss 5.410759f
C2779 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtn_1_0.RESET_B dvss 0.192338f
C2780 x2.Td_Sd.t3 dvss 0.024416f
C2781 x2.Td_Sd.t11 dvss 0.011836f
C2782 x2.Td_Sd.t16 dvss 0.016535f
C2783 x2.Td_Sd.n0 dvss 0.042092f
C2784 x2.Td_Sd.t9 dvss 0.012427f
C2785 x2.Td_Sd.t13 dvss 0.011832f
C2786 x2.Td_Sd.n1 dvss 0.047979f
C2787 x2.Td_Sd.t7 dvss 0.080224f
C2788 x2.Td_Sd.t6 dvss 0.075636f
C2789 x2.Td_Sd.n2 dvss 0.043907f
C2790 x2.Td_Sd.n3 dvss 0.175387f
C2791 x2.Td_Sd.t10 dvss 0.019447f
C2792 x2.Td_Sd.t15 dvss 0.013749f
C2793 x2.Td_Sd.n4 dvss 0.031358f
C2794 x2.delayPulse_digital_0/sky130_fd_sc_ls__dfrtp_1_0.CLK dvss 0.039715f
C2795 x2.Td_Sd.n5 dvss 0.298324f
C2796 x2.delayPulse_digital_0/sky130_fd_sc_ls__xor2_1_0.B dvss 0.018528f
C2797 x2.Td_Sd.t17 dvss 0.014531f
C2798 x2.Td_Sd.t12 dvss 0.021477f
C2799 x2.Td_Sd.n6 dvss 0.032573f
C2800 x2.Td_Sd.n7 dvss 0.015271f
C2801 x2.Td_Sd.t14 dvss 0.012886f
C2802 x2.Td_Sd.t8 dvss 0.021476f
C2803 x2.Td_Sd.n8 dvss 0.04742f
C2804 x2.Td_Sd.n9 dvss 0.226043f
C2805 x2.Td_Sd.n10 dvss 0.667997f
C2806 x2.Td_Sd.t5 dvss 0.034373f
C2807 x2.Td_Sd.t0 dvss 0.034038f
C2808 x2.Td_Sd.n11 dvss 0.295675f
C2809 x2.Td_Sd.n12 dvss 0.576755f
C2810 x2.Td_Sd.t4 dvss 0.024479f
C2811 x2.Td_Sd.t1 dvss 0.034383f
C2812 x2.Td_Sd.t2 dvss 0.034068f
C2813 x2.Td_Sd.n13 dvss 0.255204f
C2814 x2.Td_Sd.n14 dvss 0.19562f
C2815 a_35262_n291454.t3 dvss 0.013031f
C2816 a_35262_n291454.t2 dvss 0.013031f
C2817 a_35262_n291454.t4 dvss 0.013031f
C2818 a_35262_n291454.n0 dvss 0.027136f
C2819 a_35262_n291454.n1 dvss 0.020684f
C2820 a_35262_n291454.t27 dvss 0.025216f
C2821 a_35262_n291454.t21 dvss 0.027163f
C2822 a_35262_n291454.t18 dvss 0.025216f
C2823 a_35262_n291454.t12 dvss 0.027163f
C2824 a_35262_n291454.t23 dvss 0.025216f
C2825 a_35262_n291454.t15 dvss 0.027163f
C2826 a_35262_n291454.t29 dvss 0.025216f
C2827 a_35262_n291454.t24 dvss 0.036818f
C2828 a_35262_n291454.n2 dvss 0.066638f
C2829 a_35262_n291454.n3 dvss 0.04429f
C2830 a_35262_n291454.n4 dvss 0.035354f
C2831 a_35262_n291454.t11 dvss 0.025216f
C2832 a_35262_n291454.t7 dvss 0.027163f
C2833 a_35262_n291454.t25 dvss 0.025216f
C2834 a_35262_n291454.t17 dvss 0.027163f
C2835 a_35262_n291454.t6 dvss 0.025216f
C2836 a_35262_n291454.t26 dvss 0.027163f
C2837 a_35262_n291454.t16 dvss 0.025216f
C2838 a_35262_n291454.t10 dvss 0.036818f
C2839 a_35262_n291454.n5 dvss 0.066638f
C2840 a_35262_n291454.n6 dvss 0.04429f
C2841 a_35262_n291454.n7 dvss 0.035354f
C2842 a_35262_n291454.n8 dvss 0.049284f
C2843 a_35262_n291454.t20 dvss 0.010154f
C2844 a_35262_n291454.t9 dvss 0.010154f
C2845 a_35262_n291454.t13 dvss 0.010154f
C2846 a_35262_n291454.t19 dvss 0.021305f
C2847 a_35262_n291454.n9 dvss 0.060234f
C2848 a_35262_n291454.n10 dvss 0.041836f
C2849 a_35262_n291454.n11 dvss 0.0329f
C2850 a_35262_n291454.t28 dvss 0.010154f
C2851 a_35262_n291454.t14 dvss 0.010154f
C2852 a_35262_n291454.t22 dvss 0.010154f
C2853 a_35262_n291454.t8 dvss 0.021305f
C2854 a_35262_n291454.n12 dvss 0.060234f
C2855 a_35262_n291454.n13 dvss 0.041836f
C2856 a_35262_n291454.n14 dvss 0.0329f
C2857 a_35262_n291454.n15 dvss 0.049989f
C2858 a_35262_n291454.n16 dvss 0.697535f
C2859 a_35262_n291454.n17 dvss 0.277362f
C2860 a_35262_n291454.n18 dvss 0.275887f
C2861 a_35262_n291454.n19 dvss 0.026997f
C2862 a_35262_n291454.t5 dvss 0.013031f
C2863 dvdd.t107 dvss 0.016816f
C2864 dvdd.t346 dvss 0.016695f
C2865 dvdd.n0 dvss 0.158752f
C2866 dvdd.t104 dvss 0.01681f
C2867 dvdd.t105 dvss 0.016694f
C2868 dvdd.n1 dvss 0.157416f
C2869 dvdd.n2 dvss 0.010087f
C2870 dvdd.n3 dvss 0.010017f
C2871 dvdd.n4 dvss 0.088685f
C2872 dvdd.n5 dvss 0.010087f
C2873 dvdd.n6 dvss 0.010017f
C2874 dvdd.n7 dvss 0.088685f
C2875 dvdd.n8 dvss 0.010087f
C2876 dvdd.n9 dvss 0.010017f
C2877 dvdd.n10 dvss 0.088685f
C2878 dvdd.n11 dvss 0.010087f
C2879 dvdd.n12 dvss 0.010017f
C2880 dvdd.n13 dvss 0.088685f
C2881 dvdd.n14 dvss 0.010087f
C2882 dvdd.n15 dvss 0.010017f
C2883 dvdd.n16 dvss 0.088685f
C2884 dvdd.n17 dvss 0.010087f
C2885 dvdd.n18 dvss 0.010017f
C2886 dvdd.n19 dvss 0.088685f
C2887 dvdd.n20 dvss 0.010087f
C2888 dvdd.n21 dvss 0.010017f
C2889 dvdd.n22 dvss 0.088685f
C2890 dvdd.n23 dvss 0.010087f
C2891 dvdd.n24 dvss 0.010017f
C2892 dvdd.n25 dvss 0.088685f
C2893 dvdd.n26 dvss 0.010087f
C2894 dvdd.n27 dvss 0.010017f
C2895 dvdd.n28 dvss 0.088685f
C2896 dvdd.n29 dvss 0.010087f
C2897 dvdd.n30 dvss 0.010017f
C2898 dvdd.n31 dvss 0.088685f
C2899 dvdd.n32 dvss 0.010087f
C2900 dvdd.n33 dvss 0.010017f
C2901 dvdd.n34 dvss 0.088685f
C2902 dvdd.n35 dvss 0.010087f
C2903 dvdd.n36 dvss 0.010017f
C2904 dvdd.n37 dvss 0.088685f
C2905 dvdd.n38 dvss 0.010087f
C2906 dvdd.n39 dvss 0.010017f
C2907 dvdd.n40 dvss 0.088685f
C2908 dvdd.n41 dvss 0.010087f
C2909 dvdd.n42 dvss 0.010017f
C2910 dvdd.n43 dvss 0.088685f
C2911 dvdd.n44 dvss 0.010087f
C2912 dvdd.n45 dvss 0.010017f
C2913 dvdd.n46 dvss 0.088685f
C2914 dvdd.n47 dvss 0.010087f
C2915 dvdd.n48 dvss 0.010017f
C2916 dvdd.n49 dvss 0.088685f
C2917 dvdd.n50 dvss 0.010087f
C2918 dvdd.n51 dvss 0.010017f
C2919 dvdd.n52 dvss 0.088685f
C2920 dvdd.n53 dvss 0.010087f
C2921 dvdd.n54 dvss 0.010017f
C2922 dvdd.n55 dvss 0.088685f
C2923 dvdd.n56 dvss 0.010087f
C2924 dvdd.n57 dvss 0.010017f
C2925 dvdd.n58 dvss 0.088685f
C2926 dvdd.n59 dvss 0.010087f
C2927 dvdd.n60 dvss 0.010017f
C2928 dvdd.n61 dvss 0.088685f
C2929 dvdd.n62 dvss 0.010087f
C2930 dvdd.n63 dvss 0.010017f
C2931 dvdd.n64 dvss 0.088685f
C2932 dvdd.n65 dvss 0.010087f
C2933 dvdd.n66 dvss 0.010017f
C2934 dvdd.n67 dvss 0.088685f
C2935 dvdd.n68 dvss 0.010087f
C2936 dvdd.n69 dvss 0.010017f
C2937 dvdd.n70 dvss 0.088685f
C2938 dvdd.n71 dvss 0.010087f
C2939 dvdd.n72 dvss 0.010017f
C2940 dvdd.n73 dvss 0.088685f
C2941 dvdd.n74 dvss 0.010087f
C2942 dvdd.n75 dvss 0.010017f
C2943 dvdd.n76 dvss 0.088685f
C2944 dvdd.n77 dvss 0.010087f
C2945 dvdd.n78 dvss 0.010017f
C2946 dvdd.n79 dvss 0.088685f
C2947 dvdd.t139 dvss 0.016749f
C2948 dvdd.t297 dvss 0.016686f
C2949 dvdd.n80 dvss 0.092367f
C2950 dvdd.t294 dvss 0.016749f
C2951 dvdd.t266 dvss 0.016686f
C2952 dvdd.n81 dvss 0.092367f
C2953 dvdd.n82 dvss 0.503936f
C2954 dvdd.n83 dvss 0.123087f
C2955 dvdd.n84 dvss 0.123087f
C2956 dvdd.n85 dvss 0.123087f
C2957 dvdd.n86 dvss 0.123087f
C2958 dvdd.n87 dvss 0.123087f
C2959 dvdd.n88 dvss 0.123087f
C2960 dvdd.n89 dvss 0.123087f
C2961 dvdd.n90 dvss 0.123087f
C2962 dvdd.n91 dvss 0.123087f
C2963 dvdd.n92 dvss 0.123087f
C2964 dvdd.n93 dvss 0.123087f
C2965 dvdd.n94 dvss 0.123087f
C2966 dvdd.n95 dvss 0.097569f
C2967 dvdd.n96 dvss 0.229231f
C2968 dvdd.n97 dvss 0.170358f
C2969 dvdd.n98 dvss 0.161633f
C2970 dvdd.n99 dvss 0.293236f
C2971 dvdd.n100 dvss 0.293236f
C2972 dvdd.t265 dvss 0.211341f
C2973 dvdd.t292 dvss 0.139578f
C2974 dvdd.t98 dvss 0.139578f
C2975 dvdd.t38 dvss 0.139578f
C2976 dvdd.t31 dvss 0.139578f
C2977 dvdd.t162 dvss 0.139578f
C2978 dvdd.t5 dvss 0.139578f
C2979 dvdd.t45 dvss 0.139578f
C2980 dvdd.t73 dvss 0.139578f
C2981 dvdd.t268 dvss 0.139578f
C2982 dvdd.t7 dvss 0.139578f
C2983 dvdd.t100 dvss 0.139578f
C2984 dvdd.t29 dvss 0.139578f
C2985 dvdd.t303 dvss 0.211341f
C2986 dvdd.t188 dvss 0.139578f
C2987 dvdd.t186 dvss 0.139578f
C2988 dvdd.t25 dvss 0.139578f
C2989 dvdd.t21 dvss 0.139578f
C2990 dvdd.t23 dvss 0.139578f
C2991 dvdd.t192 dvss 0.139578f
C2992 dvdd.t27 dvss 0.139578f
C2993 dvdd.t77 dvss 0.139578f
C2994 dvdd.t205 dvss 0.139578f
C2995 dvdd.t311 dvss 0.139578f
C2996 dvdd.t57 dvss 0.139578f
C2997 dvdd.t47 dvss 0.139578f
C2998 dvdd.n101 dvss 0.112148f
C2999 dvdd.n102 dvss 0.120564f
C3000 dvdd.t96 dvss 0.139578f
C3001 dvdd.n103 dvss 0.120564f
C3002 dvdd.n104 dvss 0.184345f
C3003 dvdd.n105 dvss 0.498899f
C3004 dvdd.n106 dvss 0.321206f
C3005 dvdd.n107 dvss 0.091133f
C3006 dvdd.n108 dvss 0.229138f
C3007 dvdd.n109 dvss 0.184345f
C3008 dvdd.n110 dvss 0.112121f
C3009 dvdd.n111 dvss 0.120564f
C3010 dvdd.n112 dvss 0.120564f
C3011 dvdd.n113 dvss 0.161717f
C3012 dvdd.n114 dvss 0.293236f
C3013 dvdd.t138 dvss 0.211341f
C3014 dvdd.t70 dvss 0.139578f
C3015 dvdd.t255 dvss 0.139578f
C3016 dvdd.t53 dvss 0.139578f
C3017 dvdd.t259 dvss 0.139578f
C3018 dvdd.t51 dvss 0.139578f
C3019 dvdd.t270 dvss 0.139578f
C3020 dvdd.t112 dvss 0.139578f
C3021 dvdd.t146 dvss 0.139578f
C3022 dvdd.t257 dvss 0.139578f
C3023 dvdd.t79 dvss 0.139578f
C3024 dvdd.t82 dvss 0.139578f
C3025 dvdd.t195 dvss 0.139578f
C3026 dvdd.t148 dvss 0.139578f
C3027 dvdd.t84 dvss 0.139578f
C3028 dvdd.t295 dvss 0.139578f
C3029 dvdd.t227 dvss 0.139578f
C3030 dvdd.t63 dvss 0.139578f
C3031 dvdd.t94 dvss 0.139578f
C3032 dvdd.t224 dvss 0.139578f
C3033 dvdd.t92 dvss 0.139578f
C3034 dvdd.t229 dvss 0.139578f
C3035 dvdd.t231 dvss 0.139578f
C3036 dvdd.t90 dvss 0.139578f
C3037 dvdd.t280 dvss 0.139578f
C3038 dvdd.t283 dvss 0.139578f
C3039 dvdd.t200 dvss 0.211341f
C3040 dvdd.n115 dvss 0.293236f
C3041 dvdd.n116 dvss 0.170358f
C3042 dvdd.n117 dvss 0.498899f
C3043 dvdd.n118 dvss 0.321243f
C3044 dvdd.n119 dvss 0.025517f
C3045 dvdd.n120 dvss 0.031953f
C3046 dvdd.n121 dvss 0.123087f
C3047 dvdd.n122 dvss 0.123087f
C3048 dvdd.n123 dvss 0.123087f
C3049 dvdd.n124 dvss 0.123087f
C3050 dvdd.n125 dvss 0.123087f
C3051 dvdd.n126 dvss 0.123087f
C3052 dvdd.n127 dvss 0.123087f
C3053 dvdd.n128 dvss 0.123087f
C3054 dvdd.n129 dvss 0.123087f
C3055 dvdd.n130 dvss 0.123087f
C3056 dvdd.n131 dvss 0.123087f
C3057 dvdd.n132 dvss 0.123087f
C3058 dvdd.n133 dvss 0.29967f
C3059 dvdd.t118 dvss 24.4391f
C3060 dvdd.t349 dvss 39.8508f
C3061 dvdd.n134 dvss 5.13447f
C3062 dvdd.n135 dvss 0.721979f
C3063 dvdd.n136 dvss 0.785317f
C3064 dvdd.n137 dvss 0.153772f
C3065 dvdd.t20 dvss 0.016811f
C3066 dvdd.t179 dvss 0.016695f
C3067 dvdd.n138 dvss 0.150665f
C3068 dvdd.t72 dvss 0.016816f
C3069 dvdd.t18 dvss 0.016695f
C3070 dvdd.n139 dvss 0.146505f
C3071 dvdd.t178 dvss 0.015913f
C3072 dvdd.t177 dvss 0.015786f
C3073 dvdd.n140 dvss 0.149069f
C3074 dvdd.n141 dvss 0.010092f
C3075 dvdd.n142 dvss 0.01014f
C3076 dvdd.n143 dvss 0.149154f
C3077 dvdd.n144 dvss 0.015386f
C3078 dvdd.n145 dvss 0.034414f
C3079 dvdd.n146 dvss 0.022758f
C3080 dvdd.n147 dvss 0.17421f
C3081 dvdd.t308 dvss 0.127147f
C3082 dvdd.n148 dvss 0.022758f
C3083 dvdd.n149 dvss 0.033433f
C3084 dvdd.n150 dvss 0.17421f
C3085 dvdd.t59 dvss 0.146944f
C3086 dvdd.n151 dvss 0.015599f
C3087 dvdd.n152 dvss 0.196169f
C3088 dvdd.t61 dvss 0.127147f
C3089 dvdd.n153 dvss 0.023376f
C3090 dvdd.n154 dvss 0.058124f
C3091 dvdd.n155 dvss 0.023376f
C3092 dvdd.n156 dvss 0.023376f
C3093 dvdd.n157 dvss 0.022758f
C3094 dvdd.n158 dvss 0.023376f
C3095 dvdd.n159 dvss 0.023376f
C3096 dvdd.t305 dvss 0.146944f
C3097 dvdd.n160 dvss 0.058124f
C3098 dvdd.n161 dvss 0.023376f
C3099 dvdd.n162 dvss 0.176362f
C3100 dvdd.n163 dvss 0.07866f
C3101 dvdd.n164 dvss 0.273354f
C3102 dvdd.n165 dvss 0.560925f
C3103 dvdd.n166 dvss 0.198017f
C3104 dvdd.t243 dvss 0.029768f
C3105 dvdd.n167 dvss 0.045347f
C3106 dvdd.t65 dvss 0.163579f
C3107 dvdd.n168 dvss 0.015576f
C3108 dvdd.n169 dvss 0.056158f
C3109 dvdd.t2 dvss 0.021427f
C3110 dvdd.n170 dvss 0.017502f
C3111 dvdd.n171 dvss 0.023531f
C3112 dvdd.t348 dvss 0.02542f
C3113 dvdd.n172 dvss 0.018054f
C3114 dvdd.n173 dvss 0.018354f
C3115 dvdd.n174 dvss 0.02984f
C3116 dvdd.n175 dvss 0.023531f
C3117 dvdd.t241 dvss 0.01009f
C3118 dvdd.n176 dvss 0.020003f
C3119 dvdd.n177 dvss 0.01735f
C3120 dvdd.t125 dvss 0.029334f
C3121 dvdd.n178 dvss 0.036755f
C3122 dvdd.n179 dvss 0.023531f
C3123 dvdd.t161 dvss 0.017776f
C3124 dvdd.n181 dvss 0.023028f
C3125 dvdd.n182 dvss 0.023531f
C3126 dvdd.n183 dvss 0.012791f
C3127 dvdd.t109 dvss 0.0228f
C3128 dvdd.n185 dvss 0.023531f
C3129 dvdd.n186 dvss 0.014311f
C3130 dvdd.n188 dvss 0.02856f
C3131 dvdd.n189 dvss 0.023531f
C3132 dvdd.t339 dvss 0.027219f
C3133 dvdd.t286 dvss 0.022656f
C3134 dvdd.n191 dvss 0.023531f
C3135 dvdd.n193 dvss 0.026996f
C3136 dvdd.n194 dvss 0.023531f
C3137 dvdd.n195 dvss 0.022409f
C3138 dvdd.n196 dvss 0.029108f
C3139 dvdd.n197 dvss 0.017648f
C3140 dvdd.n198 dvss 0.023531f
C3141 dvdd.n199 dvss 0.023531f
C3142 dvdd.n201 dvss 0.021886f
C3143 dvdd.n202 dvss 0.016409f
C3144 dvdd.n203 dvss 0.034768f
C3145 dvdd.n204 dvss 0.023531f
C3146 dvdd.n205 dvss 0.023531f
C3147 dvdd.n206 dvss 0.023531f
C3148 dvdd.n208 dvss 0.028818f
C3149 dvdd.n211 dvss 0.023531f
C3150 dvdd.n212 dvss 0.023531f
C3151 dvdd.n213 dvss 0.023531f
C3152 dvdd.n215 dvss 0.027392f
C3153 dvdd.n216 dvss 0.040783f
C3154 dvdd.n219 dvss 0.023531f
C3155 dvdd.n220 dvss 0.023531f
C3156 dvdd.n222 dvss 0.017785f
C3157 dvdd.n225 dvss 0.023531f
C3158 dvdd.n226 dvss 0.023531f
C3159 dvdd.n227 dvss 0.023531f
C3160 dvdd.n229 dvss 0.025389f
C3161 dvdd.n231 dvss 0.017163f
C3162 dvdd.n233 dvss 0.023531f
C3163 dvdd.n234 dvss 0.023531f
C3164 dvdd.n236 dvss 0.018129f
C3165 dvdd.n238 dvss 0.023882f
C3166 dvdd.n239 dvss 0.01843f
C3167 dvdd.n241 dvss 0.017648f
C3168 dvdd.n242 dvss 0.017648f
C3169 dvdd.n243 dvss 0.023531f
C3170 dvdd.n246 dvss 0.022696f
C3171 dvdd.n247 dvss 0.024815f
C3172 dvdd.n249 dvss 0.023531f
C3173 dvdd.n250 dvss 0.023531f
C3174 dvdd.n251 dvss 0.023531f
C3175 dvdd.n254 dvss 0.023159f
C3176 dvdd.n255 dvss 0.038702f
C3177 dvdd.n257 dvss 0.017648f
C3178 dvdd.n258 dvss 0.011766f
C3179 dvdd.n259 dvss 0.024471f
C3180 dvdd.t350 dvss 0.050971f
C3181 dvdd.t1 dvss 0.021185f
C3182 dvdd.n260 dvss 0.056057f
C3183 dvdd.n261 dvss 0.015382f
C3184 dvdd.n262 dvss 0.034243f
C3185 dvdd.n264 dvss 0.025515f
C3186 dvdd.t208 dvss 0.012227f
C3187 dvdd.n265 dvss 0.122693f
C3188 dvdd.t210 dvss 0.012257f
C3189 dvdd.n266 dvss 0.215692f
C3190 dvdd.n267 dvss 0.043472f
C3191 dvdd.n268 dvss 0.033066f
C3192 dvdd.n269 dvss 0.16039f
C3193 dvdd.n270 dvss 0.16039f
C3194 dvdd.t207 dvss 0.139368f
C3195 dvdd.n271 dvss 0.030312f
C3196 dvdd.n272 dvss 0.030312f
C3197 dvdd.t209 dvss 0.139368f
C3198 dvdd.n273 dvss 0.054102f
C3199 dvdd.n274 dvss 0.030312f
C3200 dvdd.n275 dvss 0.062777f
C3201 dvdd.n276 dvss 0.096076f
C3202 dvdd.n277 dvss 0.221308f
C3203 dvdd.n278 dvss 0.011766f
C3204 dvdd.n279 dvss 0.030936f
C3205 dvdd.n280 dvss 0.076096f
C3206 dvdd.t0 dvss 0.071373f
C3207 dvdd.t248 dvss 0.067175f
C3208 dvdd.t244 dvss 0.125952f
C3209 dvdd.t246 dvss 0.100762f
C3210 dvdd.n281 dvss 0.072416f
C3211 dvdd.t128 dvss 0.033587f
C3212 dvdd.t122 dvss 0.100062f
C3213 dvdd.t347 dvss 0.069974f
C3214 dvdd.t136 dvss 0.058778f
C3215 dvdd.t35 dvss 0.062976f
C3216 dvdd.t132 dvss 0.10566f
C3217 dvdd.t130 dvss 0.111258f
C3218 dvdd.t240 dvss 0.062976f
C3219 dvdd.t126 dvss 0.07977f
C3220 dvdd.t75 dvss 0.067874f
C3221 dvdd.t134 dvss 0.069974f
C3222 dvdd.t164 dvss 0.065076f
C3223 dvdd.t124 dvss 0.081869f
C3224 dvdd.t327 dvss 0.069974f
C3225 dvdd.t325 dvss 0.060877f
C3226 dvdd.t217 dvss 0.062976f
C3227 dvdd.t171 dvss 0.065441f
C3228 dvdd.n282 dvss 0.282722f
C3229 dvdd.t160 dvss 0.067793f
C3230 dvdd.t36 dvss 0.132221f
C3231 dvdd.t212 dvss 0.076889f
C3232 dvdd.t108 dvss 0.122161f
C3233 dvdd.n283 dvss 0.581491f
C3234 dvdd.t222 dvss 0.046461f
C3235 dvdd.t111 dvss 0.062411f
C3236 dvdd.t214 dvss 0.062411f
C3237 dvdd.t66 dvss 0.054089f
C3238 dvdd.t15 dvss 0.054089f
C3239 dvdd.t203 dvss 0.085988f
C3240 dvdd.t219 dvss 0.068652f
C3241 dvdd.t169 dvss 0.063798f
C3242 dvdd.t338 dvss 0.07765f
C3243 dvdd.t211 dvss 0.056984f
C3244 dvdd.n284 dvss 1.03314f
C3245 dvdd.t223 dvss 0.103561f
C3246 dvdd.t110 dvss 0.058778f
C3247 dvdd.t67 dvss 0.058778f
C3248 dvdd.t120 dvss 0.08047f
C3249 dvdd.t215 dvss 0.075572f
C3250 dvdd.t9 dvss 0.062976f
C3251 dvdd.t250 dvss 0.062976f
C3252 dvdd.t329 dvss 0.074872f
C3253 dvdd.t252 dvss 0.135749f
C3254 dvdd.t331 dvss 0.179832f
C3255 dvdd.t242 dvss 0.070673f
C3256 dvdd.t141 dvss 0.186371f
C3257 dvdd.n285 dvss 0.222482f
C3258 dvdd.n286 dvss 0.083701f
C3259 dvdd.n287 dvss 0.78871f
C3260 dvdd.t288 dvss 0.022611f
C3261 dvdd.t290 dvss 0.022593f
C3262 dvdd.n288 dvss 0.012793f
C3263 dvdd.t302 dvss 0.022713f
C3264 dvdd.t117 dvss 0.022704f
C3265 dvdd.t44 dvss 0.022717f
C3266 dvdd.n289 dvss 0.195471f
C3267 dvdd.n290 dvss 0.049709f
C3268 dvdd.n291 dvss 0.081239f
C3269 dvdd.n292 dvss 0.028243f
C3270 dvdd.n293 dvss 0.028243f
C3271 dvdd.t43 dvss 0.333359f
C3272 dvdd.n294 dvss 0.019375f
C3273 dvdd.t151 dvss 0.333359f
C3274 dvdd.n295 dvss 0.028243f
C3275 dvdd.n296 dvss 0.028243f
C3276 dvdd.n297 dvss 0.028243f
C3277 dvdd.n298 dvss 0.017736f
C3278 dvdd.n299 dvss 0.028243f
C3279 dvdd.n300 dvss 0.028243f
C3280 dvdd.t55 dvss 0.333359f
C3281 dvdd.n301 dvss 0.019375f
C3282 dvdd.t144 dvss 0.333359f
C3283 dvdd.n302 dvss 0.028243f
C3284 dvdd.n303 dvss 0.017736f
C3285 dvdd.n304 dvss 0.081239f
C3286 dvdd.n305 dvss 0.028243f
C3287 dvdd.t184 dvss 0.333359f
C3288 dvdd.n306 dvss 0.019375f
C3289 dvdd.t40 dvss 0.333359f
C3290 dvdd.n307 dvss 0.028243f
C3291 dvdd.n308 dvss 0.017736f
C3292 dvdd.n309 dvss 0.028243f
C3293 dvdd.n310 dvss 0.028243f
C3294 dvdd.t156 dvss 0.333359f
C3295 dvdd.n311 dvss 0.019375f
C3296 dvdd.t33 dvss 0.333359f
C3297 dvdd.n312 dvss 0.028056f
C3298 dvdd.n313 dvss 0.037111f
C3299 dvdd.n314 dvss 0.017736f
C3300 dvdd.n315 dvss 0.473076f
C3301 dvdd.n316 dvss 0.017736f
C3302 dvdd.n317 dvss 0.017736f
C3303 dvdd.n318 dvss 0.037111f
C3304 dvdd.n319 dvss 0.017736f
C3305 dvdd.n320 dvss 0.473076f
C3306 dvdd.n321 dvss 0.017736f
C3307 dvdd.n322 dvss 0.017736f
C3308 dvdd.n323 dvss 0.037111f
C3309 dvdd.n324 dvss 0.017736f
C3310 dvdd.n325 dvss 0.473076f
C3311 dvdd.n326 dvss 0.017736f
C3312 dvdd.n327 dvss 0.017736f
C3313 dvdd.n328 dvss 0.017736f
C3314 dvdd.n329 dvss 0.017736f
C3315 dvdd.n330 dvss 0.037111f
C3316 dvdd.n331 dvss 0.037111f
C3317 dvdd.n332 dvss 0.037111f
C3318 dvdd.t299 dvss 0.333359f
C3319 dvdd.n333 dvss 0.017736f
C3320 dvdd.n334 dvss 0.017736f
C3321 dvdd.n335 dvss 0.473076f
C3322 dvdd.t116 dvss 0.333359f
C3323 dvdd.n336 dvss 0.019375f
C3324 dvdd.n337 dvss 0.028243f
C3325 dvdd.n338 dvss 0.017736f
C3326 dvdd.n339 dvss 0.081239f
C3327 dvdd.n340 dvss 0.028243f
C3328 dvdd.t13 dvss 0.333359f
C3329 dvdd.n341 dvss 0.019375f
C3330 dvdd.t11 dvss 0.333359f
C3331 dvdd.n342 dvss 0.028243f
C3332 dvdd.n343 dvss 0.028243f
C3333 dvdd.n344 dvss 0.017736f
C3334 dvdd.n345 dvss 0.028056f
C3335 dvdd.n346 dvss 0.028056f
C3336 dvdd.t14 dvss 0.333359f
C3337 dvdd.n347 dvss 0.019375f
C3338 dvdd.t12 dvss 0.333359f
C3339 dvdd.n348 dvss 0.026818f
C3340 dvdd.n349 dvss 0.017736f
C3341 dvdd.n350 dvss 0.02634f
C3342 dvdd.n351 dvss 0.026583f
C3343 dvdd.t320 dvss 0.07231f
C3344 dvdd.n352 dvss 0.359097f
C3345 dvdd.n353 dvss 0.017736f
C3346 dvdd.n354 dvss 0.030985f
C3347 dvdd.n355 dvss 0.020692f
C3348 dvdd.n356 dvss 0.035516f
C3349 dvdd.n357 dvss 0.037111f
C3350 dvdd.n358 dvss 0.017736f
C3351 dvdd.n359 dvss 0.473076f
C3352 dvdd.n360 dvss 0.017736f
C3353 dvdd.n361 dvss 0.017736f
C3354 dvdd.n362 dvss 0.019375f
C3355 dvdd.n363 dvss 0.037111f
C3356 dvdd.n364 dvss 0.019375f
C3357 dvdd.n365 dvss 0.030985f
C3358 dvdd.n366 dvss 0.020692f
C3359 dvdd.n367 dvss 0.026627f
C3360 dvdd.n368 dvss 0.026863f
C3361 dvdd.t287 dvss 0.07231f
C3362 dvdd.n369 dvss 0.013139f
C3363 dvdd.n370 dvss 0.012964f
C3364 dvdd.n371 dvss 0.122559f
C3365 dvdd.t317 dvss 0.161777f
C3366 dvdd.n372 dvss 0.243878f
C3367 dvdd.n373 dvss 0.139655f
C3368 dvdd.n374 dvss 0.030553f
C3369 dvdd.n375 dvss 0.035516f
C3370 dvdd.n376 dvss 0.026583f
C3371 dvdd.n377 dvss 0.026583f
C3372 dvdd.n378 dvss 0.212026f
C3373 dvdd.t289 dvss 0.161777f
C3374 dvdd.n379 dvss 0.122559f
C3375 dvdd.n380 dvss 0.026021f
C3376 dvdd.n381 dvss 0.096208f
C3377 dvdd.n382 dvss 0.075917f
C3378 dvdd.n383 dvss 0.07237f
C3379 dvdd.n384 dvss 0.019375f
C3380 dvdd.n385 dvss 0.193643f
C3381 dvdd.n386 dvss 0.028822f
C3382 dvdd.n387 dvss 0.028822f
C3383 dvdd.n388 dvss 0.028243f
C3384 dvdd.n389 dvss 0.017736f
C3385 dvdd.n390 dvss 0.473076f
C3386 dvdd.n391 dvss 0.017736f
C3387 dvdd.n392 dvss 0.017736f
C3388 dvdd.n393 dvss 0.019375f
C3389 dvdd.n394 dvss 0.028243f
C3390 dvdd.n395 dvss 0.019375f
C3391 dvdd.n396 dvss 0.019375f
C3392 dvdd.n397 dvss 0.193643f
C3393 dvdd.n398 dvss 0.019375f
C3394 dvdd.n399 dvss 0.07237f
C3395 dvdd.n400 dvss 0.081239f
C3396 dvdd.n401 dvss 0.07237f
C3397 dvdd.n402 dvss 0.019375f
C3398 dvdd.n403 dvss 0.193643f
C3399 dvdd.n404 dvss 0.019375f
C3400 dvdd.n405 dvss 0.019375f
C3401 dvdd.n406 dvss 0.037111f
C3402 dvdd.n407 dvss 0.019375f
C3403 dvdd.n408 dvss 0.037111f
C3404 dvdd.n409 dvss 0.019375f
C3405 dvdd.n410 dvss 0.037111f
C3406 dvdd.n411 dvss 0.019375f
C3407 dvdd.n412 dvss 0.037111f
C3408 dvdd.n413 dvss 0.019375f
C3409 dvdd.n414 dvss 0.028243f
C3410 dvdd.n415 dvss 0.028822f
C3411 dvdd.n416 dvss 0.028822f
C3412 dvdd.n417 dvss 0.028822f
C3413 dvdd.n418 dvss 0.037111f
C3414 dvdd.n419 dvss 0.017736f
C3415 dvdd.n420 dvss 0.017736f
C3416 dvdd.n421 dvss 0.432889f
C3417 dvdd.t262 dvss 0.173485f
C3418 dvdd.n422 dvss 0.105593f
C3419 dvdd.t154 dvss 0.201142f
C3420 dvdd.n423 dvss 0.218839f
C3421 dvdd.n424 dvss 0.038376f
C3422 dvdd.t263 dvss 0.022711f
C3423 dvdd.t34 dvss 0.022709f
C3424 dvdd.t254 dvss 0.022729f
C3425 dvdd.t41 dvss 0.022617f
C3426 dvdd.t185 dvss 0.022618f
C3427 dvdd.t145 dvss 0.022617f
C3428 dvdd.t298 dvss 0.022639f
C3429 dvdd.t166 dvss 0.022615f
C3430 dvdd.t143 dvss 0.022619f
C3431 dvdd.t165 dvss 0.022625f
C3432 dvdd.t300 dvss 0.022761f
C3433 dvdd.n425 dvss 0.342702f
C3434 dvdd.n426 dvss 0.193172f
C3435 dvdd.n427 dvss 0.193978f
C3436 dvdd.n428 dvss 0.196133f
C3437 dvdd.n429 dvss 0.195638f
C3438 dvdd.n430 dvss 0.194717f
C3439 dvdd.n431 dvss 0.186648f
C3440 dvdd.n432 dvss 0.206548f
C3441 dvdd.n433 dvss 0.19369f
C3442 dvdd.n434 dvss 0.157197f
C3443 dvdd.t155 dvss 0.022708f
C3444 dvdd.n435 dvss 0.010144f
C3445 dvdd.n436 dvss 0.010026f
C3446 dvdd.n437 dvss 0.166932f
C3447 dvdd.t4 dvss 0.015929f
C3448 dvdd.t221 dvss 0.015831f
C3449 dvdd.n438 dvss 0.184981f
C3450 dvdd.n439 dvss 0.122584f
C3451 dvdd.n440 dvss 0.080141f
C3452 dvdd.n441 dvss 0.085297f
C3453 dvdd.n442 dvss 0.027602f
C3454 dvdd.n443 dvss 0.02575f
C3455 dvdd.n444 dvss 0.319784f
C3456 dvdd.n445 dvss 0.315786f
C3457 dvdd.n446 dvss 0.027602f
C3458 dvdd.n447 dvss 0.02575f
C3459 dvdd.n448 dvss 0.042234f
C3460 dvdd.n449 dvss 0.285039f
C3461 dvdd.t273 dvss 0.237411f
C3462 dvdd.n450 dvss 0.159712f
C3463 dvdd.n451 dvss 0.030253f
C3464 dvdd.t275 dvss 0.209858f
C3465 dvdd.n452 dvss 0.095935f
C3466 dvdd.n453 dvss 0.030253f
C3467 dvdd.n454 dvss 0.030253f
C3468 dvdd.n455 dvss 0.028991f
C3469 dvdd.n456 dvss 0.028955f
C3470 dvdd.n457 dvss 0.027602f
C3471 dvdd.n458 dvss 0.028991f
C3472 dvdd.n459 dvss 0.028955f
C3473 dvdd.n460 dvss 0.02575f
C3474 dvdd.n461 dvss 0.02575f
C3475 dvdd.n462 dvss 0.011254f
C3476 dvdd.t49 dvss 0.315786f
C3477 dvdd.n463 dvss 0.02575f
C3478 dvdd.n464 dvss 0.070837f
C3479 dvdd.t182 dvss 0.01593f
C3480 dvdd.t181 dvss 0.015827f
C3481 dvdd.n465 dvss 0.184101f
C3482 dvdd.n466 dvss 0.102604f
C3483 dvdd.t50 dvss 0.01593f
C3484 dvdd.t313 dvss 0.015824f
C3485 dvdd.n467 dvss 0.182181f
C3486 dvdd.t175 dvss 0.022801f
C3487 dvdd.t316 dvss 0.022633f
C3488 dvdd.n468 dvss 0.165986f
C3489 dvdd.t336 dvss 0.022642f
C3490 dvdd.n469 dvss 0.204848f
C3491 dvdd.t322 dvss 0.022036f
C3492 dvdd.n470 dvss 0.016677f
C3493 dvdd.n471 dvss 0.079032f
C3494 dvdd.n472 dvss 0.072059f
C3495 dvdd.n473 dvss 0.072059f
C3496 dvdd.n474 dvss 0.023234f
C3497 dvdd.t324 dvss 0.022036f
C3498 dvdd.n475 dvss 0.200979f
C3499 dvdd.n476 dvss 0.375987f
C3500 dvdd.t323 dvss 0.274356f
C3501 dvdd.n477 dvss 0.131412f
C3502 dvdd.t321 dvss 0.274356f
C3503 dvdd.n478 dvss 0.375987f
C3504 dvdd.n479 dvss 0.023437f
C3505 dvdd.n480 dvss 0.156204f
C3506 dvdd.n481 dvss 0.216075f
C3507 dvdd.n483 dvss 3.69214f
C3508 dvdd.n484 dvss 2.51047f
C3509 dvdd.t337 dvss 0.02263f
C3510 dvdd.n485 dvss 0.259791f
C3511 dvdd.n486 dvss 0.252671f
C3512 dvdd.n487 dvss 0.127262f
C3513 dvdd.n488 dvss 0.171057f
C3514 dvdd.n489 dvss 0.091558f
C3515 dvdd.n490 dvss 0.026622f
C3516 dvdd.n491 dvss 0.026622f
C3517 dvdd.n492 dvss 0.034921f
C3518 dvdd.t174 dvss 0.345766f
C3519 dvdd.n493 dvss 0.029839f
C3520 dvdd.n494 dvss 0.105017f
C3521 dvdd.n495 dvss 0.028248f
C3522 dvdd.n496 dvss 0.033229f
C3523 dvdd.n497 dvss 0.044097f
C3524 dvdd.n498 dvss 0.028955f
C3525 dvdd.n499 dvss 0.302152f
C3526 dvdd.t335 dvss 0.368667f
C3527 dvdd.n501 dvss 0.027649f
C3528 dvdd.n502 dvss 0.028955f
C3529 dvdd.n503 dvss 0.029819f
C3530 dvdd.n504 dvss 0.029839f
C3531 dvdd.n505 dvss 0.028955f
C3532 dvdd.n506 dvss 0.033265f
C3533 dvdd.n507 dvss 0.396029f
C3534 dvdd.n508 dvss 0.105017f
C3535 dvdd.n509 dvss 0.064454f
C3536 dvdd.n510 dvss 0.049941f
C3537 dvdd.n511 dvss 0.043345f
C3538 dvdd.n512 dvss 0.061087f
C3539 dvdd.n513 dvss 0.029043f
C3540 dvdd.n514 dvss 0.018874f
C3541 dvdd.n515 dvss 0.010726f
C3542 dvdd.n516 dvss 0.046242f
C3543 dvdd.n517 dvss 0.278811f
C3544 dvdd.n518 dvss 0.263821f
C3545 dvdd.n519 dvss 0.040923f
C3546 dvdd.n520 dvss 0.026622f
C3547 dvdd.n521 dvss 0.04573f
C3548 dvdd.n522 dvss 0.085297f
C3549 dvdd.n523 dvss 0.028955f
C3550 dvdd.n524 dvss 0.028991f
C3551 dvdd.n525 dvss 0.315786f
C3552 dvdd.t180 dvss 0.315786f
C3553 dvdd.n526 dvss 0.011254f
C3554 dvdd.n527 dvss 0.011254f
C3555 dvdd.n528 dvss 0.02575f
C3556 dvdd.n529 dvss 0.011254f
C3557 dvdd.n530 dvss 0.011254f
C3558 dvdd.t3 dvss 0.315786f
C3559 dvdd.n531 dvss 0.011254f
C3560 dvdd.n532 dvss 0.052231f
C3561 dvdd.n533 dvss 0.169603f
C3562 dvdd.n534 dvss 0.407286f
C3563 dvdd.n535 dvss 0.328458f
C3564 dvdd.t272 dvss 0.022874f
C3565 dvdd.t157 dvss 0.02287f
C3566 dvdd.t86 dvss 0.022869f
C3567 dvdd.t279 dvss 0.022864f
C3568 dvdd.t267 dvss 0.022859f
C3569 dvdd.t56 dvss 0.022869f
C3570 dvdd.t152 dvss 0.022702f
C3571 dvdd.n536 dvss 0.234296f
C3572 dvdd.n537 dvss 0.253464f
C3573 dvdd.n538 dvss 0.249293f
C3574 dvdd.n539 dvss 0.250198f
C3575 dvdd.n540 dvss 0.249565f
C3576 dvdd.n541 dvss 0.24591f
C3577 dvdd.n542 dvss 0.348111f
C3578 dvdd.n543 dvss 0.578068f
C3579 dvdd.n544 dvss 0.212113f
C3580 dvdd.n545 dvss 0.197734f
C3581 dvdd.n546 dvss 0.118825f
C3582 dvdd.n547 dvss 0.039334f
C3583 dvdd.n548 dvss 0.110729f
C3584 dvdd.n549 dvss 0.028822f
C3585 dvdd.n550 dvss 0.193643f
C3586 dvdd.n551 dvss 0.019375f
C3587 dvdd.n552 dvss 0.019375f
C3588 dvdd.n553 dvss 0.028243f
C3589 dvdd.n554 dvss 0.019375f
C3590 dvdd.n555 dvss 0.019375f
C3591 dvdd.n556 dvss 0.193643f
C3592 dvdd.n557 dvss 0.019375f
C3593 dvdd.n558 dvss 0.07237f
C3594 dvdd.n559 dvss 0.081239f
C3595 dvdd.n560 dvss 0.07237f
C3596 dvdd.n561 dvss 0.019375f
C3597 dvdd.n562 dvss 0.193643f
C3598 dvdd.n563 dvss 0.019375f
C3599 dvdd.n564 dvss 0.019375f
C3600 dvdd.n565 dvss 0.028243f
C3601 dvdd.n566 dvss 0.019375f
C3602 dvdd.n567 dvss 0.019375f
C3603 dvdd.n568 dvss 0.193643f
C3604 dvdd.n569 dvss 0.019375f
C3605 dvdd.n570 dvss 0.067713f
C3606 dvdd.n571 dvss 0.329976f
C3607 dvdd.n572 dvss 0.732514f
C3608 dvdd.n573 dvss 0.219039f
C3609 dvdd.n574 dvss 0.297843f
C3610 dvdd.n575 dvss 0.471964f
C3611 dvdd.n576 dvss 0.489275f
C3612 dvdd.n577 dvss 0.253761f
C3613 dvdd.n578 dvss 0.976776f
C3614 dvdd.n579 dvss 0.590627f
C3615 dvdd.n580 dvss 0.20887f
C3616 dvdd.n581 dvss 0.09561f
C3617 dvdd.n582 dvss 0.095832f
C3618 dvdd.n583 dvss 0.029454f
C3619 dvdd.n584 dvss 0.027602f
C3620 dvdd.t19 dvss 0.209858f
C3621 dvdd.n585 dvss 0.014958f
C3622 dvdd.t176 dvss 0.343543f
C3623 dvdd.n586 dvss 0.027602f
C3624 dvdd.n587 dvss 0.028991f
C3625 dvdd.n588 dvss 0.041932f
C3626 dvdd.n589 dvss 0.285039f
C3627 dvdd.n590 dvss 0.029454f
C3628 dvdd.t103 dvss 0.237411f
C3629 dvdd.n591 dvss 0.028991f
C3630 dvdd.n592 dvss 0.323781f
C3631 dvdd.t106 dvss 0.209858f
C3632 dvdd.n593 dvss 0.153564f
C3633 dvdd.n594 dvss 0.030253f
C3634 dvdd.n595 dvss 0.095935f
C3635 dvdd.n596 dvss 0.030253f
C3636 dvdd.n597 dvss 0.030253f
C3637 dvdd.n598 dvss 0.029454f
C3638 dvdd.n599 dvss 0.014958f
C3639 dvdd.n600 dvss 0.038286f
C3640 dvdd.n601 dvss 0.122703f
C3641 dvdd.n602 dvss 0.026622f
C3642 dvdd.n603 dvss 0.276987f
C3643 dvdd.n605 dvss 0.026622f
C3644 dvdd.n606 dvss 0.026622f
C3645 dvdd.n607 dvss 0.027602f
C3646 dvdd.n608 dvss 0.028991f
C3647 dvdd.n609 dvss 0.028991f
C3648 dvdd.n610 dvss 0.319784f
C3649 dvdd.t17 dvss 0.209858f
C3650 dvdd.n611 dvss 0.095935f
C3651 dvdd.n612 dvss 0.014958f
C3652 dvdd.n613 dvss 0.058128f
C3653 dvdd.n614 dvss 0.210785f
C3654 dvdd.n615 dvss 0.454222f
C3655 dvdd.n616 dvss 0.071168f
C3656 x2.VT2.t2 dvss 1.46595f
C3657 x2.VT2.n0 dvss 0.012889f
C3658 x2.VT2.t1 dvss 2.35105f
C3659 x2.VT2.t0 dvss 2.7556f
C3660 x2.VT2.n2 dvss 0.233308f
C3661 x2.VT2.t3 dvss 1.3743f
.ends

