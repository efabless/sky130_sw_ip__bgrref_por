magic
tech sky130A
magscale 1 2
timestamp 1731360119
<< isosubstrate >>
rect 3992 -292617 17571 -279609
<< nwell >>
rect 3668 -279490 17889 -279310
rect 3668 -292646 3908 -279490
rect 17460 -279508 17889 -279490
rect 17709 -285270 17889 -279508
rect 32362 -283550 38526 -283370
rect 32362 -285270 32542 -283550
rect 17709 -285450 32542 -285270
rect 38286 -286171 38526 -283550
rect 38152 -287265 38526 -286171
rect 38286 -292646 38526 -287265
rect 3668 -292890 38526 -292646
<< mvpsubdiff >>
rect 3489 -279177 3549 -279143
rect 17991 -279177 18056 -279143
rect 3489 -279203 3523 -279177
rect 18022 -279198 18056 -279177
rect 18022 -285103 18056 -285071
rect 32195 -283237 32255 -283203
rect 38627 -283237 38687 -283203
rect 32195 -283263 32229 -283237
rect 38653 -283263 38687 -283237
rect 32195 -285103 32229 -285078
rect 18022 -285137 18081 -285103
rect 32163 -285137 32229 -285103
rect 3489 -293013 3523 -292987
rect 38653 -293013 38687 -292987
rect 3489 -293047 3549 -293013
rect 38627 -293047 38687 -293013
<< mvnsubdiff >>
rect 3734 -279410 3794 -279376
rect 17759 -279410 17823 -279376
rect 3734 -279436 3768 -279410
rect 17789 -279441 17823 -279410
rect 32428 -283470 32488 -283436
rect 38400 -283470 38460 -283436
rect 32428 -283496 32462 -283470
rect 17789 -285336 17823 -285296
rect 32428 -285336 32462 -285302
rect 17789 -285370 17857 -285336
rect 32388 -285370 32462 -285336
rect 38426 -283496 38460 -283470
rect 3734 -292790 3768 -292764
rect 38426 -292790 38460 -292764
rect 3734 -292824 3794 -292790
rect 38400 -292824 38460 -292790
<< mvpsubdiffcont >>
rect 3549 -279177 17991 -279143
rect 3489 -292987 3523 -279203
rect 18022 -285071 18056 -279198
rect 32255 -283237 38627 -283203
rect 32195 -285078 32229 -283263
rect 18081 -285137 32163 -285103
rect 38653 -292987 38687 -283263
rect 3549 -293047 38627 -293013
<< mvnsubdiffcont >>
rect 3794 -279410 17759 -279376
rect 3734 -292764 3768 -279436
rect 17789 -285296 17823 -279441
rect 32488 -283470 38400 -283436
rect 32428 -285302 32462 -283496
rect 17857 -285370 32388 -285336
rect 38426 -292764 38460 -283496
rect 3794 -292824 38400 -292790
<< locali >>
rect 3489 -279177 3549 -279143
rect 17991 -279177 18056 -279143
rect 3489 -279198 18056 -279177
rect 3489 -279203 18022 -279198
rect 3523 -279214 18022 -279203
rect 3523 -279260 3551 -279214
rect 3523 -279310 17939 -279260
rect 3523 -279347 3633 -279310
rect 3523 -292843 3540 -279347
rect 3583 -292843 3633 -279347
rect 3734 -279410 3794 -279376
rect 17759 -279410 17823 -279376
rect 3734 -279436 17823 -279410
rect 3768 -279441 17823 -279436
rect 3768 -279446 17789 -279441
rect 3768 -279490 3804 -279446
rect 3768 -279530 17709 -279490
rect 3768 -279548 3895 -279530
rect 3768 -292656 3802 -279548
rect 3844 -292656 3895 -279548
rect 7353 -279717 15350 -279714
rect 7292 -279760 15350 -279717
rect 7292 -279801 7498 -279760
rect 7292 -289021 7360 -279801
rect 7412 -279816 7498 -279801
rect 15275 -279816 15350 -279760
rect 7412 -279903 15350 -279816
rect 7412 -288909 7481 -279903
rect 11766 -280590 12544 -279903
rect 11766 -288849 12025 -280590
rect 12322 -288849 12544 -280590
rect 11766 -288909 12544 -288849
rect 15161 -279905 15350 -279903
rect 15161 -288182 15216 -279905
rect 15268 -287795 15350 -279905
rect 17669 -285450 17709 -279530
rect 17753 -285296 17789 -279446
rect 17889 -285220 17939 -279310
rect 17985 -285071 18022 -279214
rect 17985 -285103 18056 -285071
rect 32195 -283237 32255 -283203
rect 38627 -283237 38687 -283203
rect 32195 -283263 38687 -283237
rect 32229 -283274 38653 -283263
rect 32229 -283320 32257 -283274
rect 38510 -283306 38653 -283274
rect 38510 -283320 38595 -283306
rect 32229 -283370 38595 -283320
rect 32229 -283407 32362 -283370
rect 32229 -285078 32266 -283407
rect 32195 -285103 32266 -285078
rect 17985 -285137 18081 -285103
rect 32163 -285137 32266 -285103
rect 17985 -285174 32266 -285137
rect 32312 -285220 32362 -283407
rect 17889 -285270 32362 -285220
rect 32428 -283470 32488 -283436
rect 38400 -283470 38460 -283436
rect 32428 -283496 38460 -283470
rect 17753 -285336 17823 -285296
rect 32462 -283506 38426 -283496
rect 32462 -283550 32498 -283506
rect 38319 -283525 38426 -283506
rect 38319 -283550 38363 -283525
rect 32462 -283590 38363 -283550
rect 32462 -283608 32582 -283590
rect 32462 -285302 32498 -283608
rect 32428 -285336 32498 -285302
rect 17753 -285370 17857 -285336
rect 32388 -285370 32498 -285336
rect 17753 -285406 32498 -285370
rect 32542 -285450 32582 -283608
rect 17669 -285490 32582 -285450
rect 15928 -287795 16180 -287790
rect 15268 -287903 16180 -287795
rect 15268 -288182 15414 -287903
rect 15161 -288909 15414 -288182
rect 15928 -287906 16180 -287903
rect 15928 -288909 16024 -287906
rect 7412 -288987 16024 -288909
rect 7412 -289021 7479 -288987
rect 7292 -289047 7479 -289021
rect 9970 -289013 16024 -288987
rect 9970 -289047 13305 -289013
rect 7292 -289062 13305 -289047
rect 15607 -289046 16024 -289013
rect 16160 -289046 16180 -287906
rect 15607 -289062 16180 -289046
rect 7292 -289065 16180 -289062
rect 7292 -289098 11061 -289065
rect 11030 -289118 11061 -289098
rect 13220 -289098 16180 -289065
rect 13220 -289118 13244 -289098
rect 11030 -289355 13244 -289118
rect 3768 -292692 3895 -292656
rect 38324 -292692 38363 -283590
rect 3768 -292732 38363 -292692
rect 3768 -292764 3821 -292732
rect 3734 -292769 3821 -292764
rect 38284 -292746 38363 -292732
rect 38402 -292746 38426 -283525
rect 38284 -292764 38426 -292746
rect 38284 -292769 38460 -292764
rect 3734 -292790 38460 -292769
rect 3734 -292824 3794 -292790
rect 38400 -292824 38460 -292790
rect 3523 -292877 3633 -292843
rect 38553 -292873 38595 -283370
rect 38634 -292873 38653 -283306
rect 38553 -292877 38653 -292873
rect 3523 -292942 38653 -292877
rect 3523 -292981 3593 -292942
rect 38616 -292981 38653 -292942
rect 3523 -292987 38653 -292981
rect 3489 -293013 38687 -292987
rect 3489 -293047 3549 -293013
rect 38627 -293047 38687 -293013
<< viali >>
rect 3551 -279260 17985 -279214
rect 3540 -292843 3583 -279347
rect 3804 -279490 17753 -279446
rect 3802 -292656 3844 -279548
rect 7360 -289021 7412 -279801
rect 7498 -279816 15275 -279760
rect 15216 -288182 15268 -279905
rect 17709 -285406 17753 -279490
rect 17939 -285174 17985 -279260
rect 32257 -283320 38510 -283274
rect 32266 -285174 32312 -283407
rect 17939 -285220 32312 -285174
rect 32498 -283550 38319 -283506
rect 32498 -285406 32542 -283608
rect 17709 -285450 32542 -285406
rect 7479 -289047 9970 -288987
rect 13305 -289062 15607 -289013
rect 16024 -289046 16160 -287906
rect 11061 -289118 13220 -289065
rect 3821 -292769 38284 -292732
rect 38363 -292746 38402 -283525
rect 38595 -292873 38634 -283306
rect 3593 -292981 38616 -292942
<< metal1 >>
rect 3493 -279214 18049 -279150
rect 3493 -279260 3551 -279214
rect 3493 -279302 17939 -279260
rect 3502 -279347 3612 -279302
rect 3502 -292843 3540 -279347
rect 3583 -292843 3612 -279347
rect 3756 -279436 17806 -279393
rect 3756 -279446 6368 -279436
rect 3756 -279490 3804 -279446
rect 3756 -279508 6368 -279490
rect 17754 -279508 17806 -279436
rect 3756 -279519 17709 -279508
rect 3756 -279548 3877 -279519
rect 3756 -289178 3802 -279548
rect 3844 -289178 3877 -279548
rect 7295 -279715 7513 -279713
rect 7295 -279760 15350 -279715
rect 7295 -279801 7498 -279760
rect 7295 -279840 7360 -279801
rect 7412 -279816 7498 -279801
rect 15275 -279816 15350 -279760
rect 7295 -288899 7327 -279840
rect 7412 -279894 15350 -279816
rect 7412 -279997 7513 -279894
rect 15145 -279905 15350 -279894
rect 7412 -280429 7676 -279997
rect 7772 -280429 8008 -279997
rect 8104 -280429 8340 -279997
rect 8436 -280429 8672 -279997
rect 8768 -280429 9004 -279997
rect 9100 -280429 9336 -279997
rect 9432 -280429 9668 -279997
rect 9764 -280429 10000 -279997
rect 10096 -280429 10332 -279997
rect 10428 -280429 10664 -279997
rect 10760 -280429 10996 -279997
rect 11092 -280429 11328 -279997
rect 11424 -280429 11660 -279997
rect 12125 -280116 12716 -280115
rect 12124 -280429 12716 -280116
rect 12800 -280429 13038 -279996
rect 13134 -280429 13372 -279996
rect 13468 -280429 13706 -279996
rect 13802 -280429 14040 -279996
rect 14136 -280429 14374 -279996
rect 14470 -280429 14708 -279996
rect 14804 -280429 15042 -279996
rect 7295 -289021 7360 -288899
rect 7412 -288907 7513 -280429
rect 12124 -281147 12198 -280429
rect 7606 -288829 7842 -288397
rect 7938 -288829 8174 -288397
rect 8270 -288829 8506 -288397
rect 8602 -288829 8838 -288397
rect 8934 -288829 9170 -288397
rect 9266 -288829 9502 -288397
rect 9598 -288829 9834 -288397
rect 9930 -288829 10166 -288397
rect 10262 -288829 10498 -288397
rect 10594 -288829 10830 -288397
rect 10926 -288829 11162 -288397
rect 11258 -288829 11494 -288397
rect 11588 -288747 12197 -288397
rect 11827 -288868 11874 -288747
rect 7412 -288976 10050 -288907
rect 7412 -289021 7467 -288976
rect 7295 -289052 7467 -289021
rect 10015 -289052 10050 -288976
rect 7295 -289094 10050 -289052
rect 10468 -288915 11874 -288868
rect 7901 -289096 8874 -289094
rect 3756 -289467 3772 -289178
rect 3870 -289467 3877 -289178
rect 10468 -289262 10515 -288915
rect 12407 -288953 12455 -280429
rect 15145 -288182 15216 -279905
rect 15268 -288182 15350 -279905
rect 17680 -285450 17709 -279519
rect 17753 -285353 17806 -279508
rect 17897 -285220 17939 -279302
rect 17985 -285110 18049 -279214
rect 32199 -283274 38674 -283210
rect 32199 -283320 32257 -283274
rect 38510 -283306 38674 -283274
rect 38510 -283320 38595 -283306
rect 32199 -283362 38595 -283320
rect 32202 -283407 32354 -283362
rect 32202 -285110 32266 -283407
rect 17985 -285174 32266 -285110
rect 32312 -285220 32354 -283407
rect 17897 -285262 32354 -285220
rect 32445 -283457 38440 -283453
rect 32445 -283506 38447 -283457
rect 32445 -283550 32498 -283506
rect 38319 -283525 38447 -283506
rect 38319 -283550 38363 -283525
rect 32445 -283579 38363 -283550
rect 32445 -283608 32571 -283579
rect 32445 -285353 32498 -283608
rect 17753 -285406 32498 -285353
rect 32542 -285450 32571 -283608
rect 17680 -285479 32571 -285450
rect 15145 -288235 15350 -288182
rect 15415 -287747 16312 -287471
rect 16605 -287747 16614 -287471
rect 15415 -288324 15543 -287747
rect 15648 -288025 15692 -287747
rect 16006 -287906 16180 -287786
rect 15579 -288067 15746 -288025
rect 15648 -288340 15692 -288067
rect 15579 -288382 15746 -288340
rect 12634 -288829 12872 -288396
rect 12968 -288829 13206 -288396
rect 13302 -288829 13540 -288396
rect 13636 -288829 13874 -288396
rect 13970 -288829 14208 -288396
rect 14304 -288829 14542 -288396
rect 14638 -288829 14876 -288396
rect 14983 -288829 15545 -288394
rect 15648 -288448 15692 -288382
rect 15579 -288490 15746 -288448
rect 15648 -288762 15692 -288490
rect 15579 -288829 15746 -288762
rect 15791 -288763 15952 -288074
rect 10784 -289001 12455 -288953
rect 13056 -288976 15663 -288972
rect 10784 -289210 10832 -289001
rect 13056 -289013 13403 -288976
rect 15496 -289013 15663 -288976
rect 13056 -289043 13305 -289013
rect 11027 -289062 13305 -289043
rect 15607 -289062 15663 -289013
rect 11027 -289065 15663 -289062
rect 11027 -289118 11061 -289065
rect 13220 -289092 15663 -289065
rect 16006 -289046 16024 -287906
rect 16160 -289046 16180 -287906
rect 13220 -289118 13240 -289092
rect 16006 -289102 16180 -289046
rect 11027 -289355 13240 -289118
rect 3756 -292656 3802 -289467
rect 3844 -292656 3877 -289467
rect 17538 -290701 17586 -289045
rect 16990 -290749 17586 -290701
rect 3986 -292610 17746 -292563
rect 3986 -292611 23772 -292610
rect 3756 -292703 3877 -292656
rect 38334 -292703 38363 -283579
rect 3756 -292732 38363 -292703
rect 3756 -292769 3821 -292732
rect 38284 -292746 38363 -292732
rect 38402 -292746 38447 -283525
rect 38284 -292769 38447 -292746
rect 3756 -292802 38447 -292769
rect 3756 -292805 38380 -292802
rect 3758 -292809 38380 -292805
rect 3502 -292902 3612 -292843
rect 38562 -292873 38595 -283362
rect 38634 -283362 38674 -283306
rect 38634 -292873 38672 -283362
rect 38562 -292902 38672 -292873
rect 3502 -292927 38672 -292902
rect 3502 -292942 17403 -292927
rect 24818 -292942 38672 -292927
rect 3502 -292981 3593 -292942
rect 38616 -292981 38672 -292942
rect 3502 -293001 17403 -292981
rect 24818 -293001 38672 -292981
rect 3502 -293032 38672 -293001
rect 38562 -293043 38672 -293032
<< via1 >>
rect 6368 -279446 17754 -279436
rect 6368 -279490 17753 -279446
rect 6368 -279508 17709 -279490
rect 17709 -279508 17753 -279490
rect 17753 -279508 17754 -279446
rect 7327 -288899 7360 -279840
rect 7360 -288899 7403 -279840
rect 7467 -288987 10015 -288976
rect 7467 -289047 7479 -288987
rect 7479 -289047 9970 -288987
rect 9970 -289047 10015 -288987
rect 7467 -289052 10015 -289047
rect 3772 -289467 3802 -289178
rect 3802 -289467 3844 -289178
rect 3844 -289467 3870 -289178
rect 16312 -287747 16605 -287471
rect 13403 -289013 15496 -288976
rect 13403 -289041 15496 -289013
rect 16024 -289046 16160 -287906
rect 16786 -289428 17380 -289293
rect 5791 -292476 9241 -292342
rect 12676 -292483 16558 -292395
rect 17403 -292942 24818 -292927
rect 17403 -292981 24818 -292942
rect 17403 -293001 24818 -292981
<< metal2 >>
rect 6314 -279436 17834 -279397
rect 6314 -279497 6368 -279436
rect 6312 -279508 6368 -279497
rect 17754 -279508 17834 -279436
rect 6312 -279652 17834 -279508
rect 6312 -279660 6605 -279652
rect 7200 -279840 7466 -279763
rect 7200 -288899 7327 -279840
rect 7403 -288806 7466 -279840
rect 16312 -284876 16605 -279652
rect 39229 -284155 39429 -284118
rect 37892 -284274 39429 -284155
rect 39229 -284318 39429 -284274
rect 24237 -284876 24891 -284875
rect 16312 -285327 24891 -284876
rect 39229 -284905 39429 -284868
rect 37892 -285024 39429 -284905
rect 39229 -285068 39429 -285024
rect 16312 -287471 16605 -285327
rect 24237 -285850 24891 -285327
rect 24238 -286408 24891 -285850
rect 15937 -287906 16181 -287878
rect 15937 -288806 16024 -287906
rect 7403 -288899 16024 -288806
rect 7200 -288976 16024 -288899
rect 7200 -289052 7467 -288976
rect 10015 -289041 13403 -288976
rect 15496 -289041 16024 -288976
rect 10015 -289046 16024 -289041
rect 16160 -289046 16181 -287906
rect 10015 -289052 16181 -289046
rect 7200 -289070 16181 -289052
rect 7200 -289072 16078 -289070
rect 3464 -289178 4428 -289169
rect 3464 -289467 3772 -289178
rect 3870 -289467 4428 -289178
rect 16312 -289183 16605 -287747
rect 3464 -289479 4428 -289467
rect 15582 -289476 16605 -289183
rect 16747 -288187 17828 -287923
rect 16747 -289293 17438 -288187
rect 39296 -289256 39496 -289188
rect 16747 -289428 16786 -289293
rect 17380 -289428 17438 -289293
rect 38044 -289340 39496 -289256
rect 39296 -289388 39496 -289340
rect 16747 -289466 17438 -289428
rect 35038 -290006 39195 -290005
rect 35038 -290381 39497 -290006
rect 39301 -290786 39501 -290729
rect 37952 -290871 39501 -290786
rect 37952 -291076 38037 -290871
rect 39301 -290929 39501 -290871
rect 4462 -292342 9298 -292313
rect 3569 -292649 4341 -292449
rect 4462 -292476 5791 -292342
rect 9241 -292476 9298 -292342
rect 4462 -292805 9298 -292476
rect 12630 -292395 16597 -292360
rect 12630 -292483 12676 -292395
rect 16558 -292483 16597 -292395
rect 12630 -292805 16597 -292483
rect 4462 -292806 16600 -292805
rect 3564 -293345 16600 -292806
rect 4462 -293347 16600 -293345
rect 17324 -292927 17872 -292805
rect 17324 -293001 17403 -292927
rect 17324 -293003 17872 -293001
rect 17324 -293338 24877 -293003
rect 17324 -293347 17872 -293338
<< metal3 >>
rect 32079 -284981 32641 -284194
<< metal4 >>
rect 32079 -284981 32641 -284194
<< metal5 >>
rect 32079 -284981 32641 -284194
use por_via_4cut  por_via_4cut_3
timestamp 1718283729
transform -1 0 20299 0 -1 -300491
box 15948 -7932 16222 -7868
use por_via_4cut  por_via_4cut_18
timestamp 1718283729
transform 0 -1 9676 1 0 -305162
box 15948 -7932 16222 -7868
use sky130_fd_pr__res_xhigh_po_0p35_MNWQZD  R12 paramcells
timestamp 1731359787
transform 1 0 13835 0 1 -284412
box -1363 -4582 1363 4582
use sky130_fd_pr__res_xhigh_po_0p35_WGPHGK  R1 paramcells
timestamp 1731359787
transform 1 0 9633 0 1 -284414
box -2193 -4582 2193 4582
use sky130_fd_pr__res_xhigh_po_0p35_YTHETB  R10 paramcells
timestamp 1731359787
transform 1 0 12163 0 1 -284732
box -201 -4182 201 4182
use comparator_final  x1
timestamp 1731357245
transform 1 0 6296 0 1 -286728
box -1988 -5804 11208 -1484
use delayPulse_final  x2
timestamp 1731360119
transform 1 0 1048 0 1 -2959
box 1311 -297437 38614 -274935
use sky130_fd_pr__nfet_05v0_nvt_CZFQWY  XM2 paramcells
timestamp 1726591550
transform 1 0 15668 0 1 -288416
box -318 -567 318 567
<< labels >>
flabel metal2 39296 -289388 39496 -289188 0 FreeSans 256 0 0 0 porb
port 5 nsew
flabel metal2 39301 -290929 39501 -290729 0 FreeSans 256 0 0 0 por
port 1 nsew
flabel metal2 24555 -293294 24755 -293094 0 FreeSans 256 0 0 0 dvss
port 6 nsew
flabel metal2 39292 -290256 39492 -290056 0 FreeSans 256 0 0 0 dvdd
port 4 nsew
flabel metal2 3491 -289455 3691 -289255 0 FreeSans 256 0 0 0 avdd
port 3 nsew
flabel metal2 3569 -292649 3769 -292449 0 FreeSans 256 0 0 0 vbg
port 0 nsew
flabel metal2 3612 -293264 3812 -293064 0 FreeSans 256 0 0 0 avss
port 2 nsew
flabel metal2 39229 -285068 39429 -284868 0 FreeSans 256 0 0 0 porb_h[1]
port 8 nsew
flabel metal2 39229 -284318 39429 -284118 0 FreeSans 256 0 0 0 porb_h[0]
port 7 nsew
<< end >>
